magic
tech sky130A
magscale 1 2
timestamp 1755207335
<< viali >>
rect 2605 21641 2639 21675
rect 11713 21641 11747 21675
rect 20269 21641 20303 21675
rect 2881 21505 2915 21539
rect 11621 21505 11655 21539
rect 20085 21505 20119 21539
rect 22385 20009 22419 20043
rect 22201 19805 22235 19839
rect 4261 18921 4295 18955
rect 10977 18921 11011 18955
rect 4445 18717 4479 18751
rect 10793 18717 10827 18751
rect 4261 18377 4295 18411
rect 10885 18377 10919 18411
rect 19165 18377 19199 18411
rect 4445 18309 4479 18343
rect 10701 18309 10735 18343
rect 1501 18241 1535 18275
rect 18981 18241 19015 18275
rect 10333 18173 10367 18207
rect 4813 18105 4847 18139
rect 1777 18037 1811 18071
rect 4445 18037 4479 18071
rect 10701 18037 10735 18071
rect 17601 17833 17635 17867
rect 18153 17833 18187 17867
rect 18337 17833 18371 17867
rect 17509 17765 17543 17799
rect 17601 17629 17635 17663
rect 17785 17629 17819 17663
rect 17325 17561 17359 17595
rect 18153 17493 18187 17527
rect 19073 10761 19107 10795
rect 18889 10625 18923 10659
rect 22201 10625 22235 10659
rect 22385 10421 22419 10455
rect 18153 10217 18187 10251
rect 18337 10217 18371 10251
rect 17969 9945 18003 9979
rect 18174 9877 18208 9911
rect 4169 8993 4203 9027
rect 4077 8925 4111 8959
rect 4261 8925 4295 8959
rect 1409 8857 1443 8891
rect 1777 8857 1811 8891
rect 3893 8857 3927 8891
rect 16773 5185 16807 5219
rect 16865 5185 16899 5219
rect 16957 5117 16991 5151
rect 17141 4981 17175 5015
rect 8217 4097 8251 4131
rect 8309 4097 8343 4131
rect 8125 4029 8159 4063
rect 8493 3893 8527 3927
rect 1777 2601 1811 2635
rect 22109 2601 22143 2635
rect 9045 2397 9079 2431
rect 16957 2397 16991 2431
rect 1501 2329 1535 2363
rect 22385 2329 22419 2363
rect 9137 2261 9171 2295
rect 17049 2261 17083 2295
<< metal1 >>
rect 1104 21786 22816 21808
rect 1104 21734 4324 21786
rect 4376 21734 4388 21786
rect 4440 21734 4452 21786
rect 4504 21734 4516 21786
rect 4568 21734 4580 21786
rect 4632 21734 9752 21786
rect 9804 21734 9816 21786
rect 9868 21734 9880 21786
rect 9932 21734 9944 21786
rect 9996 21734 10008 21786
rect 10060 21734 15180 21786
rect 15232 21734 15244 21786
rect 15296 21734 15308 21786
rect 15360 21734 15372 21786
rect 15424 21734 15436 21786
rect 15488 21734 20608 21786
rect 20660 21734 20672 21786
rect 20724 21734 20736 21786
rect 20788 21734 20800 21786
rect 20852 21734 20864 21786
rect 20916 21734 22816 21786
rect 1104 21712 22816 21734
rect 2590 21632 2596 21684
rect 2648 21632 2654 21684
rect 11146 21632 11152 21684
rect 11204 21672 11210 21684
rect 11701 21675 11759 21681
rect 11701 21672 11713 21675
rect 11204 21644 11713 21672
rect 11204 21632 11210 21644
rect 11701 21641 11713 21644
rect 11747 21641 11759 21675
rect 11701 21635 11759 21641
rect 20254 21632 20260 21684
rect 20312 21632 20318 21684
rect 2869 21539 2927 21545
rect 2869 21505 2881 21539
rect 2915 21536 2927 21539
rect 4246 21536 4252 21548
rect 2915 21508 4252 21536
rect 2915 21505 2927 21508
rect 2869 21499 2927 21505
rect 4246 21496 4252 21508
rect 4304 21496 4310 21548
rect 10962 21496 10968 21548
rect 11020 21536 11026 21548
rect 11609 21539 11667 21545
rect 11609 21536 11621 21539
rect 11020 21508 11621 21536
rect 11020 21496 11026 21508
rect 11609 21505 11621 21508
rect 11655 21505 11667 21539
rect 11609 21499 11667 21505
rect 18046 21496 18052 21548
rect 18104 21536 18110 21548
rect 20073 21539 20131 21545
rect 20073 21536 20085 21539
rect 18104 21508 20085 21536
rect 18104 21496 18110 21508
rect 20073 21505 20085 21508
rect 20119 21505 20131 21539
rect 20073 21499 20131 21505
rect 1104 21242 22816 21264
rect 1104 21190 3664 21242
rect 3716 21190 3728 21242
rect 3780 21190 3792 21242
rect 3844 21190 3856 21242
rect 3908 21190 3920 21242
rect 3972 21190 9092 21242
rect 9144 21190 9156 21242
rect 9208 21190 9220 21242
rect 9272 21190 9284 21242
rect 9336 21190 9348 21242
rect 9400 21190 14520 21242
rect 14572 21190 14584 21242
rect 14636 21190 14648 21242
rect 14700 21190 14712 21242
rect 14764 21190 14776 21242
rect 14828 21190 19948 21242
rect 20000 21190 20012 21242
rect 20064 21190 20076 21242
rect 20128 21190 20140 21242
rect 20192 21190 20204 21242
rect 20256 21190 22816 21242
rect 1104 21168 22816 21190
rect 1104 20698 22816 20720
rect 1104 20646 4324 20698
rect 4376 20646 4388 20698
rect 4440 20646 4452 20698
rect 4504 20646 4516 20698
rect 4568 20646 4580 20698
rect 4632 20646 9752 20698
rect 9804 20646 9816 20698
rect 9868 20646 9880 20698
rect 9932 20646 9944 20698
rect 9996 20646 10008 20698
rect 10060 20646 15180 20698
rect 15232 20646 15244 20698
rect 15296 20646 15308 20698
rect 15360 20646 15372 20698
rect 15424 20646 15436 20698
rect 15488 20646 20608 20698
rect 20660 20646 20672 20698
rect 20724 20646 20736 20698
rect 20788 20646 20800 20698
rect 20852 20646 20864 20698
rect 20916 20646 22816 20698
rect 1104 20624 22816 20646
rect 1104 20154 22816 20176
rect 1104 20102 3664 20154
rect 3716 20102 3728 20154
rect 3780 20102 3792 20154
rect 3844 20102 3856 20154
rect 3908 20102 3920 20154
rect 3972 20102 9092 20154
rect 9144 20102 9156 20154
rect 9208 20102 9220 20154
rect 9272 20102 9284 20154
rect 9336 20102 9348 20154
rect 9400 20102 14520 20154
rect 14572 20102 14584 20154
rect 14636 20102 14648 20154
rect 14700 20102 14712 20154
rect 14764 20102 14776 20154
rect 14828 20102 19948 20154
rect 20000 20102 20012 20154
rect 20064 20102 20076 20154
rect 20128 20102 20140 20154
rect 20192 20102 20204 20154
rect 20256 20102 22816 20154
rect 1104 20080 22816 20102
rect 22373 20043 22431 20049
rect 22373 20009 22385 20043
rect 22419 20040 22431 20043
rect 22419 20012 22876 20040
rect 22419 20009 22431 20012
rect 22373 20003 22431 20009
rect 22848 19984 22876 20012
rect 22830 19932 22836 19984
rect 22888 19932 22894 19984
rect 22186 19796 22192 19848
rect 22244 19796 22250 19848
rect 1104 19610 22816 19632
rect 1104 19558 4324 19610
rect 4376 19558 4388 19610
rect 4440 19558 4452 19610
rect 4504 19558 4516 19610
rect 4568 19558 4580 19610
rect 4632 19558 9752 19610
rect 9804 19558 9816 19610
rect 9868 19558 9880 19610
rect 9932 19558 9944 19610
rect 9996 19558 10008 19610
rect 10060 19558 15180 19610
rect 15232 19558 15244 19610
rect 15296 19558 15308 19610
rect 15360 19558 15372 19610
rect 15424 19558 15436 19610
rect 15488 19558 20608 19610
rect 20660 19558 20672 19610
rect 20724 19558 20736 19610
rect 20788 19558 20800 19610
rect 20852 19558 20864 19610
rect 20916 19558 22816 19610
rect 1104 19536 22816 19558
rect 1104 19066 22816 19088
rect 1104 19014 3664 19066
rect 3716 19014 3728 19066
rect 3780 19014 3792 19066
rect 3844 19014 3856 19066
rect 3908 19014 3920 19066
rect 3972 19014 9092 19066
rect 9144 19014 9156 19066
rect 9208 19014 9220 19066
rect 9272 19014 9284 19066
rect 9336 19014 9348 19066
rect 9400 19014 14520 19066
rect 14572 19014 14584 19066
rect 14636 19014 14648 19066
rect 14700 19014 14712 19066
rect 14764 19014 14776 19066
rect 14828 19014 19948 19066
rect 20000 19014 20012 19066
rect 20064 19014 20076 19066
rect 20128 19014 20140 19066
rect 20192 19014 20204 19066
rect 20256 19014 22816 19066
rect 1104 18992 22816 19014
rect 4246 18912 4252 18964
rect 4304 18912 4310 18964
rect 10962 18912 10968 18964
rect 11020 18912 11026 18964
rect 4246 18708 4252 18760
rect 4304 18748 4310 18760
rect 4433 18751 4491 18757
rect 4433 18748 4445 18751
rect 4304 18720 4445 18748
rect 4304 18708 4310 18720
rect 4433 18717 4445 18720
rect 4479 18717 4491 18751
rect 4433 18711 4491 18717
rect 10778 18708 10784 18760
rect 10836 18708 10842 18760
rect 1104 18522 22816 18544
rect 1104 18470 4324 18522
rect 4376 18470 4388 18522
rect 4440 18470 4452 18522
rect 4504 18470 4516 18522
rect 4568 18470 4580 18522
rect 4632 18470 9752 18522
rect 9804 18470 9816 18522
rect 9868 18470 9880 18522
rect 9932 18470 9944 18522
rect 9996 18470 10008 18522
rect 10060 18470 15180 18522
rect 15232 18470 15244 18522
rect 15296 18470 15308 18522
rect 15360 18470 15372 18522
rect 15424 18470 15436 18522
rect 15488 18470 20608 18522
rect 20660 18470 20672 18522
rect 20724 18470 20736 18522
rect 20788 18470 20800 18522
rect 20852 18470 20864 18522
rect 20916 18470 22816 18522
rect 1104 18448 22816 18470
rect 4246 18368 4252 18420
rect 4304 18368 4310 18420
rect 10778 18368 10784 18420
rect 10836 18408 10842 18420
rect 10873 18411 10931 18417
rect 10873 18408 10885 18411
rect 10836 18380 10885 18408
rect 10836 18368 10842 18380
rect 10873 18377 10885 18380
rect 10919 18377 10931 18411
rect 10873 18371 10931 18377
rect 19153 18411 19211 18417
rect 19153 18377 19165 18411
rect 19199 18408 19211 18411
rect 22186 18408 22192 18420
rect 19199 18380 22192 18408
rect 19199 18377 19211 18380
rect 19153 18371 19211 18377
rect 22186 18368 22192 18380
rect 22244 18368 22250 18420
rect 4154 18300 4160 18352
rect 4212 18340 4218 18352
rect 4433 18343 4491 18349
rect 4433 18340 4445 18343
rect 4212 18312 4445 18340
rect 4212 18300 4218 18312
rect 4433 18309 4445 18312
rect 4479 18340 4491 18343
rect 10689 18343 10747 18349
rect 10689 18340 10701 18343
rect 4479 18312 10701 18340
rect 4479 18309 4491 18312
rect 4433 18303 4491 18309
rect 10689 18309 10701 18312
rect 10735 18309 10747 18343
rect 10689 18303 10747 18309
rect 1486 18232 1492 18284
rect 1544 18232 1550 18284
rect 18966 18232 18972 18284
rect 19024 18232 19030 18284
rect 10321 18207 10379 18213
rect 10321 18204 10333 18207
rect 4448 18176 10333 18204
rect 1765 18071 1823 18077
rect 1765 18037 1777 18071
rect 1811 18068 1823 18071
rect 4062 18068 4068 18080
rect 1811 18040 4068 18068
rect 1811 18037 1823 18040
rect 1765 18031 1823 18037
rect 4062 18028 4068 18040
rect 4120 18068 4126 18080
rect 4448 18077 4476 18176
rect 10321 18173 10333 18176
rect 10367 18204 10379 18207
rect 10367 18176 15240 18204
rect 10367 18173 10379 18176
rect 10321 18167 10379 18173
rect 15212 18148 15240 18176
rect 4801 18139 4859 18145
rect 4801 18105 4813 18139
rect 4847 18105 4859 18139
rect 4801 18099 4859 18105
rect 4433 18071 4491 18077
rect 4433 18068 4445 18071
rect 4120 18040 4445 18068
rect 4120 18028 4126 18040
rect 4433 18037 4445 18040
rect 4479 18037 4491 18071
rect 4816 18068 4844 18099
rect 15194 18096 15200 18148
rect 15252 18096 15258 18148
rect 10689 18071 10747 18077
rect 10689 18068 10701 18071
rect 4816 18040 10701 18068
rect 4433 18031 4491 18037
rect 10689 18037 10701 18040
rect 10735 18068 10747 18071
rect 17494 18068 17500 18080
rect 10735 18040 17500 18068
rect 10735 18037 10747 18040
rect 10689 18031 10747 18037
rect 17494 18028 17500 18040
rect 17552 18028 17558 18080
rect 1104 17978 22816 18000
rect 1104 17926 3664 17978
rect 3716 17926 3728 17978
rect 3780 17926 3792 17978
rect 3844 17926 3856 17978
rect 3908 17926 3920 17978
rect 3972 17926 9092 17978
rect 9144 17926 9156 17978
rect 9208 17926 9220 17978
rect 9272 17926 9284 17978
rect 9336 17926 9348 17978
rect 9400 17926 14520 17978
rect 14572 17926 14584 17978
rect 14636 17926 14648 17978
rect 14700 17926 14712 17978
rect 14764 17926 14776 17978
rect 14828 17926 19948 17978
rect 20000 17926 20012 17978
rect 20064 17926 20076 17978
rect 20128 17926 20140 17978
rect 20192 17926 20204 17978
rect 20256 17926 22816 17978
rect 1104 17904 22816 17926
rect 17589 17867 17647 17873
rect 17589 17833 17601 17867
rect 17635 17864 17647 17867
rect 18046 17864 18052 17876
rect 17635 17836 18052 17864
rect 17635 17833 17647 17836
rect 17589 17827 17647 17833
rect 18046 17824 18052 17836
rect 18104 17824 18110 17876
rect 18138 17824 18144 17876
rect 18196 17824 18202 17876
rect 18325 17867 18383 17873
rect 18325 17833 18337 17867
rect 18371 17864 18383 17867
rect 18966 17864 18972 17876
rect 18371 17836 18972 17864
rect 18371 17833 18383 17836
rect 18325 17827 18383 17833
rect 18966 17824 18972 17836
rect 19024 17824 19030 17876
rect 17494 17756 17500 17808
rect 17552 17796 17558 17808
rect 18156 17796 18184 17824
rect 17552 17768 18184 17796
rect 17552 17756 17558 17768
rect 15194 17688 15200 17740
rect 15252 17728 15258 17740
rect 15252 17700 18184 17728
rect 15252 17688 15258 17700
rect 17604 17669 17632 17700
rect 17589 17663 17647 17669
rect 17589 17629 17601 17663
rect 17635 17629 17647 17663
rect 17589 17623 17647 17629
rect 17770 17620 17776 17672
rect 17828 17620 17834 17672
rect 17313 17595 17371 17601
rect 17313 17561 17325 17595
rect 17359 17592 17371 17595
rect 17788 17592 17816 17620
rect 17359 17564 17816 17592
rect 17359 17561 17371 17564
rect 17313 17555 17371 17561
rect 18156 17533 18184 17700
rect 18141 17527 18199 17533
rect 18141 17493 18153 17527
rect 18187 17524 18199 17527
rect 18230 17524 18236 17536
rect 18187 17496 18236 17524
rect 18187 17493 18199 17496
rect 18141 17487 18199 17493
rect 18230 17484 18236 17496
rect 18288 17484 18294 17536
rect 1104 17434 22816 17456
rect 1104 17382 4324 17434
rect 4376 17382 4388 17434
rect 4440 17382 4452 17434
rect 4504 17382 4516 17434
rect 4568 17382 4580 17434
rect 4632 17382 9752 17434
rect 9804 17382 9816 17434
rect 9868 17382 9880 17434
rect 9932 17382 9944 17434
rect 9996 17382 10008 17434
rect 10060 17382 15180 17434
rect 15232 17382 15244 17434
rect 15296 17382 15308 17434
rect 15360 17382 15372 17434
rect 15424 17382 15436 17434
rect 15488 17382 20608 17434
rect 20660 17382 20672 17434
rect 20724 17382 20736 17434
rect 20788 17382 20800 17434
rect 20852 17382 20864 17434
rect 20916 17382 22816 17434
rect 1104 17360 22816 17382
rect 1104 16890 22816 16912
rect 1104 16838 3664 16890
rect 3716 16838 3728 16890
rect 3780 16838 3792 16890
rect 3844 16838 3856 16890
rect 3908 16838 3920 16890
rect 3972 16838 9092 16890
rect 9144 16838 9156 16890
rect 9208 16838 9220 16890
rect 9272 16838 9284 16890
rect 9336 16838 9348 16890
rect 9400 16838 14520 16890
rect 14572 16838 14584 16890
rect 14636 16838 14648 16890
rect 14700 16838 14712 16890
rect 14764 16838 14776 16890
rect 14828 16838 19948 16890
rect 20000 16838 20012 16890
rect 20064 16838 20076 16890
rect 20128 16838 20140 16890
rect 20192 16838 20204 16890
rect 20256 16838 22816 16890
rect 1104 16816 22816 16838
rect 1104 16346 22816 16368
rect 1104 16294 4324 16346
rect 4376 16294 4388 16346
rect 4440 16294 4452 16346
rect 4504 16294 4516 16346
rect 4568 16294 4580 16346
rect 4632 16294 9752 16346
rect 9804 16294 9816 16346
rect 9868 16294 9880 16346
rect 9932 16294 9944 16346
rect 9996 16294 10008 16346
rect 10060 16294 15180 16346
rect 15232 16294 15244 16346
rect 15296 16294 15308 16346
rect 15360 16294 15372 16346
rect 15424 16294 15436 16346
rect 15488 16294 20608 16346
rect 20660 16294 20672 16346
rect 20724 16294 20736 16346
rect 20788 16294 20800 16346
rect 20852 16294 20864 16346
rect 20916 16294 22816 16346
rect 1104 16272 22816 16294
rect 1104 15802 22816 15824
rect 1104 15750 3664 15802
rect 3716 15750 3728 15802
rect 3780 15750 3792 15802
rect 3844 15750 3856 15802
rect 3908 15750 3920 15802
rect 3972 15750 9092 15802
rect 9144 15750 9156 15802
rect 9208 15750 9220 15802
rect 9272 15750 9284 15802
rect 9336 15750 9348 15802
rect 9400 15750 14520 15802
rect 14572 15750 14584 15802
rect 14636 15750 14648 15802
rect 14700 15750 14712 15802
rect 14764 15750 14776 15802
rect 14828 15750 19948 15802
rect 20000 15750 20012 15802
rect 20064 15750 20076 15802
rect 20128 15750 20140 15802
rect 20192 15750 20204 15802
rect 20256 15750 22816 15802
rect 1104 15728 22816 15750
rect 1104 15258 22816 15280
rect 1104 15206 4324 15258
rect 4376 15206 4388 15258
rect 4440 15206 4452 15258
rect 4504 15206 4516 15258
rect 4568 15206 4580 15258
rect 4632 15206 9752 15258
rect 9804 15206 9816 15258
rect 9868 15206 9880 15258
rect 9932 15206 9944 15258
rect 9996 15206 10008 15258
rect 10060 15206 15180 15258
rect 15232 15206 15244 15258
rect 15296 15206 15308 15258
rect 15360 15206 15372 15258
rect 15424 15206 15436 15258
rect 15488 15206 20608 15258
rect 20660 15206 20672 15258
rect 20724 15206 20736 15258
rect 20788 15206 20800 15258
rect 20852 15206 20864 15258
rect 20916 15206 22816 15258
rect 1104 15184 22816 15206
rect 1104 14714 22816 14736
rect 1104 14662 3664 14714
rect 3716 14662 3728 14714
rect 3780 14662 3792 14714
rect 3844 14662 3856 14714
rect 3908 14662 3920 14714
rect 3972 14662 9092 14714
rect 9144 14662 9156 14714
rect 9208 14662 9220 14714
rect 9272 14662 9284 14714
rect 9336 14662 9348 14714
rect 9400 14662 14520 14714
rect 14572 14662 14584 14714
rect 14636 14662 14648 14714
rect 14700 14662 14712 14714
rect 14764 14662 14776 14714
rect 14828 14662 19948 14714
rect 20000 14662 20012 14714
rect 20064 14662 20076 14714
rect 20128 14662 20140 14714
rect 20192 14662 20204 14714
rect 20256 14662 22816 14714
rect 1104 14640 22816 14662
rect 1104 14170 22816 14192
rect 1104 14118 4324 14170
rect 4376 14118 4388 14170
rect 4440 14118 4452 14170
rect 4504 14118 4516 14170
rect 4568 14118 4580 14170
rect 4632 14118 9752 14170
rect 9804 14118 9816 14170
rect 9868 14118 9880 14170
rect 9932 14118 9944 14170
rect 9996 14118 10008 14170
rect 10060 14118 15180 14170
rect 15232 14118 15244 14170
rect 15296 14118 15308 14170
rect 15360 14118 15372 14170
rect 15424 14118 15436 14170
rect 15488 14118 20608 14170
rect 20660 14118 20672 14170
rect 20724 14118 20736 14170
rect 20788 14118 20800 14170
rect 20852 14118 20864 14170
rect 20916 14118 22816 14170
rect 1104 14096 22816 14118
rect 1104 13626 22816 13648
rect 1104 13574 3664 13626
rect 3716 13574 3728 13626
rect 3780 13574 3792 13626
rect 3844 13574 3856 13626
rect 3908 13574 3920 13626
rect 3972 13574 9092 13626
rect 9144 13574 9156 13626
rect 9208 13574 9220 13626
rect 9272 13574 9284 13626
rect 9336 13574 9348 13626
rect 9400 13574 14520 13626
rect 14572 13574 14584 13626
rect 14636 13574 14648 13626
rect 14700 13574 14712 13626
rect 14764 13574 14776 13626
rect 14828 13574 19948 13626
rect 20000 13574 20012 13626
rect 20064 13574 20076 13626
rect 20128 13574 20140 13626
rect 20192 13574 20204 13626
rect 20256 13574 22816 13626
rect 1104 13552 22816 13574
rect 1104 13082 22816 13104
rect 1104 13030 4324 13082
rect 4376 13030 4388 13082
rect 4440 13030 4452 13082
rect 4504 13030 4516 13082
rect 4568 13030 4580 13082
rect 4632 13030 9752 13082
rect 9804 13030 9816 13082
rect 9868 13030 9880 13082
rect 9932 13030 9944 13082
rect 9996 13030 10008 13082
rect 10060 13030 15180 13082
rect 15232 13030 15244 13082
rect 15296 13030 15308 13082
rect 15360 13030 15372 13082
rect 15424 13030 15436 13082
rect 15488 13030 20608 13082
rect 20660 13030 20672 13082
rect 20724 13030 20736 13082
rect 20788 13030 20800 13082
rect 20852 13030 20864 13082
rect 20916 13030 22816 13082
rect 1104 13008 22816 13030
rect 1104 12538 22816 12560
rect 1104 12486 3664 12538
rect 3716 12486 3728 12538
rect 3780 12486 3792 12538
rect 3844 12486 3856 12538
rect 3908 12486 3920 12538
rect 3972 12486 9092 12538
rect 9144 12486 9156 12538
rect 9208 12486 9220 12538
rect 9272 12486 9284 12538
rect 9336 12486 9348 12538
rect 9400 12486 14520 12538
rect 14572 12486 14584 12538
rect 14636 12486 14648 12538
rect 14700 12486 14712 12538
rect 14764 12486 14776 12538
rect 14828 12486 19948 12538
rect 20000 12486 20012 12538
rect 20064 12486 20076 12538
rect 20128 12486 20140 12538
rect 20192 12486 20204 12538
rect 20256 12486 22816 12538
rect 1104 12464 22816 12486
rect 1104 11994 22816 12016
rect 1104 11942 4324 11994
rect 4376 11942 4388 11994
rect 4440 11942 4452 11994
rect 4504 11942 4516 11994
rect 4568 11942 4580 11994
rect 4632 11942 9752 11994
rect 9804 11942 9816 11994
rect 9868 11942 9880 11994
rect 9932 11942 9944 11994
rect 9996 11942 10008 11994
rect 10060 11942 15180 11994
rect 15232 11942 15244 11994
rect 15296 11942 15308 11994
rect 15360 11942 15372 11994
rect 15424 11942 15436 11994
rect 15488 11942 20608 11994
rect 20660 11942 20672 11994
rect 20724 11942 20736 11994
rect 20788 11942 20800 11994
rect 20852 11942 20864 11994
rect 20916 11942 22816 11994
rect 1104 11920 22816 11942
rect 1104 11450 22816 11472
rect 1104 11398 3664 11450
rect 3716 11398 3728 11450
rect 3780 11398 3792 11450
rect 3844 11398 3856 11450
rect 3908 11398 3920 11450
rect 3972 11398 9092 11450
rect 9144 11398 9156 11450
rect 9208 11398 9220 11450
rect 9272 11398 9284 11450
rect 9336 11398 9348 11450
rect 9400 11398 14520 11450
rect 14572 11398 14584 11450
rect 14636 11398 14648 11450
rect 14700 11398 14712 11450
rect 14764 11398 14776 11450
rect 14828 11398 19948 11450
rect 20000 11398 20012 11450
rect 20064 11398 20076 11450
rect 20128 11398 20140 11450
rect 20192 11398 20204 11450
rect 20256 11398 22816 11450
rect 1104 11376 22816 11398
rect 1104 10906 22816 10928
rect 1104 10854 4324 10906
rect 4376 10854 4388 10906
rect 4440 10854 4452 10906
rect 4504 10854 4516 10906
rect 4568 10854 4580 10906
rect 4632 10854 9752 10906
rect 9804 10854 9816 10906
rect 9868 10854 9880 10906
rect 9932 10854 9944 10906
rect 9996 10854 10008 10906
rect 10060 10854 15180 10906
rect 15232 10854 15244 10906
rect 15296 10854 15308 10906
rect 15360 10854 15372 10906
rect 15424 10854 15436 10906
rect 15488 10854 20608 10906
rect 20660 10854 20672 10906
rect 20724 10854 20736 10906
rect 20788 10854 20800 10906
rect 20852 10854 20864 10906
rect 20916 10854 22816 10906
rect 1104 10832 22816 10854
rect 19061 10795 19119 10801
rect 19061 10761 19073 10795
rect 19107 10761 19119 10795
rect 19061 10755 19119 10761
rect 18874 10616 18880 10668
rect 18932 10616 18938 10668
rect 19076 10656 19104 10755
rect 22189 10659 22247 10665
rect 22189 10656 22201 10659
rect 19076 10628 22201 10656
rect 22189 10625 22201 10628
rect 22235 10625 22247 10659
rect 22189 10619 22247 10625
rect 22370 10412 22376 10464
rect 22428 10412 22434 10464
rect 1104 10362 22816 10384
rect 1104 10310 3664 10362
rect 3716 10310 3728 10362
rect 3780 10310 3792 10362
rect 3844 10310 3856 10362
rect 3908 10310 3920 10362
rect 3972 10310 9092 10362
rect 9144 10310 9156 10362
rect 9208 10310 9220 10362
rect 9272 10310 9284 10362
rect 9336 10310 9348 10362
rect 9400 10310 14520 10362
rect 14572 10310 14584 10362
rect 14636 10310 14648 10362
rect 14700 10310 14712 10362
rect 14764 10310 14776 10362
rect 14828 10310 19948 10362
rect 20000 10310 20012 10362
rect 20064 10310 20076 10362
rect 20128 10310 20140 10362
rect 20192 10310 20204 10362
rect 20256 10310 22816 10362
rect 1104 10288 22816 10310
rect 18138 10208 18144 10260
rect 18196 10208 18202 10260
rect 18325 10251 18383 10257
rect 18325 10217 18337 10251
rect 18371 10248 18383 10251
rect 18874 10248 18880 10260
rect 18371 10220 18880 10248
rect 18371 10217 18383 10220
rect 18325 10211 18383 10217
rect 18874 10208 18880 10220
rect 18932 10208 18938 10260
rect 18230 10004 18236 10056
rect 18288 10004 18294 10056
rect 16850 9936 16856 9988
rect 16908 9976 16914 9988
rect 17770 9976 17776 9988
rect 16908 9948 17776 9976
rect 16908 9936 16914 9948
rect 17770 9936 17776 9948
rect 17828 9976 17834 9988
rect 17957 9979 18015 9985
rect 17957 9976 17969 9979
rect 17828 9948 17969 9976
rect 17828 9936 17834 9948
rect 17957 9945 17969 9948
rect 18003 9945 18015 9979
rect 17957 9939 18015 9945
rect 18162 9911 18220 9917
rect 18162 9877 18174 9911
rect 18208 9908 18220 9911
rect 18248 9908 18276 10004
rect 18208 9880 18276 9908
rect 18208 9877 18220 9880
rect 18162 9871 18220 9877
rect 1104 9818 22816 9840
rect 1104 9766 4324 9818
rect 4376 9766 4388 9818
rect 4440 9766 4452 9818
rect 4504 9766 4516 9818
rect 4568 9766 4580 9818
rect 4632 9766 9752 9818
rect 9804 9766 9816 9818
rect 9868 9766 9880 9818
rect 9932 9766 9944 9818
rect 9996 9766 10008 9818
rect 10060 9766 15180 9818
rect 15232 9766 15244 9818
rect 15296 9766 15308 9818
rect 15360 9766 15372 9818
rect 15424 9766 15436 9818
rect 15488 9766 20608 9818
rect 20660 9766 20672 9818
rect 20724 9766 20736 9818
rect 20788 9766 20800 9818
rect 20852 9766 20864 9818
rect 20916 9766 22816 9818
rect 1104 9744 22816 9766
rect 1104 9274 22816 9296
rect 1104 9222 3664 9274
rect 3716 9222 3728 9274
rect 3780 9222 3792 9274
rect 3844 9222 3856 9274
rect 3908 9222 3920 9274
rect 3972 9222 9092 9274
rect 9144 9222 9156 9274
rect 9208 9222 9220 9274
rect 9272 9222 9284 9274
rect 9336 9222 9348 9274
rect 9400 9222 14520 9274
rect 14572 9222 14584 9274
rect 14636 9222 14648 9274
rect 14700 9222 14712 9274
rect 14764 9222 14776 9274
rect 14828 9222 19948 9274
rect 20000 9222 20012 9274
rect 20064 9222 20076 9274
rect 20128 9222 20140 9274
rect 20192 9222 20204 9274
rect 20256 9222 22816 9274
rect 1104 9200 22816 9222
rect 4154 8984 4160 9036
rect 4212 9024 4218 9036
rect 4706 9024 4712 9036
rect 4212 8996 4712 9024
rect 4212 8984 4218 8996
rect 4706 8984 4712 8996
rect 4764 8984 4770 9036
rect 4062 8916 4068 8968
rect 4120 8916 4126 8968
rect 4249 8959 4307 8965
rect 4249 8925 4261 8959
rect 4295 8956 4307 8959
rect 8018 8956 8024 8968
rect 4295 8928 8024 8956
rect 4295 8925 4307 8928
rect 4249 8919 4307 8925
rect 8018 8916 8024 8928
rect 8076 8916 8082 8968
rect 934 8848 940 8900
rect 992 8888 998 8900
rect 1397 8891 1455 8897
rect 1397 8888 1409 8891
rect 992 8860 1409 8888
rect 992 8848 998 8860
rect 1397 8857 1409 8860
rect 1443 8857 1455 8891
rect 1397 8851 1455 8857
rect 1765 8891 1823 8897
rect 1765 8857 1777 8891
rect 1811 8888 1823 8891
rect 3881 8891 3939 8897
rect 3881 8888 3893 8891
rect 1811 8860 3893 8888
rect 1811 8857 1823 8860
rect 1765 8851 1823 8857
rect 3881 8857 3893 8860
rect 3927 8857 3939 8891
rect 3881 8851 3939 8857
rect 1104 8730 22816 8752
rect 1104 8678 4324 8730
rect 4376 8678 4388 8730
rect 4440 8678 4452 8730
rect 4504 8678 4516 8730
rect 4568 8678 4580 8730
rect 4632 8678 9752 8730
rect 9804 8678 9816 8730
rect 9868 8678 9880 8730
rect 9932 8678 9944 8730
rect 9996 8678 10008 8730
rect 10060 8678 15180 8730
rect 15232 8678 15244 8730
rect 15296 8678 15308 8730
rect 15360 8678 15372 8730
rect 15424 8678 15436 8730
rect 15488 8678 20608 8730
rect 20660 8678 20672 8730
rect 20724 8678 20736 8730
rect 20788 8678 20800 8730
rect 20852 8678 20864 8730
rect 20916 8678 22816 8730
rect 1104 8656 22816 8678
rect 1104 8186 22816 8208
rect 1104 8134 3664 8186
rect 3716 8134 3728 8186
rect 3780 8134 3792 8186
rect 3844 8134 3856 8186
rect 3908 8134 3920 8186
rect 3972 8134 9092 8186
rect 9144 8134 9156 8186
rect 9208 8134 9220 8186
rect 9272 8134 9284 8186
rect 9336 8134 9348 8186
rect 9400 8134 14520 8186
rect 14572 8134 14584 8186
rect 14636 8134 14648 8186
rect 14700 8134 14712 8186
rect 14764 8134 14776 8186
rect 14828 8134 19948 8186
rect 20000 8134 20012 8186
rect 20064 8134 20076 8186
rect 20128 8134 20140 8186
rect 20192 8134 20204 8186
rect 20256 8134 22816 8186
rect 1104 8112 22816 8134
rect 1104 7642 22816 7664
rect 1104 7590 4324 7642
rect 4376 7590 4388 7642
rect 4440 7590 4452 7642
rect 4504 7590 4516 7642
rect 4568 7590 4580 7642
rect 4632 7590 9752 7642
rect 9804 7590 9816 7642
rect 9868 7590 9880 7642
rect 9932 7590 9944 7642
rect 9996 7590 10008 7642
rect 10060 7590 15180 7642
rect 15232 7590 15244 7642
rect 15296 7590 15308 7642
rect 15360 7590 15372 7642
rect 15424 7590 15436 7642
rect 15488 7590 20608 7642
rect 20660 7590 20672 7642
rect 20724 7590 20736 7642
rect 20788 7590 20800 7642
rect 20852 7590 20864 7642
rect 20916 7590 22816 7642
rect 1104 7568 22816 7590
rect 1104 7098 22816 7120
rect 1104 7046 3664 7098
rect 3716 7046 3728 7098
rect 3780 7046 3792 7098
rect 3844 7046 3856 7098
rect 3908 7046 3920 7098
rect 3972 7046 9092 7098
rect 9144 7046 9156 7098
rect 9208 7046 9220 7098
rect 9272 7046 9284 7098
rect 9336 7046 9348 7098
rect 9400 7046 14520 7098
rect 14572 7046 14584 7098
rect 14636 7046 14648 7098
rect 14700 7046 14712 7098
rect 14764 7046 14776 7098
rect 14828 7046 19948 7098
rect 20000 7046 20012 7098
rect 20064 7046 20076 7098
rect 20128 7046 20140 7098
rect 20192 7046 20204 7098
rect 20256 7046 22816 7098
rect 1104 7024 22816 7046
rect 1104 6554 22816 6576
rect 1104 6502 4324 6554
rect 4376 6502 4388 6554
rect 4440 6502 4452 6554
rect 4504 6502 4516 6554
rect 4568 6502 4580 6554
rect 4632 6502 9752 6554
rect 9804 6502 9816 6554
rect 9868 6502 9880 6554
rect 9932 6502 9944 6554
rect 9996 6502 10008 6554
rect 10060 6502 15180 6554
rect 15232 6502 15244 6554
rect 15296 6502 15308 6554
rect 15360 6502 15372 6554
rect 15424 6502 15436 6554
rect 15488 6502 20608 6554
rect 20660 6502 20672 6554
rect 20724 6502 20736 6554
rect 20788 6502 20800 6554
rect 20852 6502 20864 6554
rect 20916 6502 22816 6554
rect 1104 6480 22816 6502
rect 1104 6010 22816 6032
rect 1104 5958 3664 6010
rect 3716 5958 3728 6010
rect 3780 5958 3792 6010
rect 3844 5958 3856 6010
rect 3908 5958 3920 6010
rect 3972 5958 9092 6010
rect 9144 5958 9156 6010
rect 9208 5958 9220 6010
rect 9272 5958 9284 6010
rect 9336 5958 9348 6010
rect 9400 5958 14520 6010
rect 14572 5958 14584 6010
rect 14636 5958 14648 6010
rect 14700 5958 14712 6010
rect 14764 5958 14776 6010
rect 14828 5958 19948 6010
rect 20000 5958 20012 6010
rect 20064 5958 20076 6010
rect 20128 5958 20140 6010
rect 20192 5958 20204 6010
rect 20256 5958 22816 6010
rect 1104 5936 22816 5958
rect 1104 5466 22816 5488
rect 1104 5414 4324 5466
rect 4376 5414 4388 5466
rect 4440 5414 4452 5466
rect 4504 5414 4516 5466
rect 4568 5414 4580 5466
rect 4632 5414 9752 5466
rect 9804 5414 9816 5466
rect 9868 5414 9880 5466
rect 9932 5414 9944 5466
rect 9996 5414 10008 5466
rect 10060 5414 15180 5466
rect 15232 5414 15244 5466
rect 15296 5414 15308 5466
rect 15360 5414 15372 5466
rect 15424 5414 15436 5466
rect 15488 5414 20608 5466
rect 20660 5414 20672 5466
rect 20724 5414 20736 5466
rect 20788 5414 20800 5466
rect 20852 5414 20864 5466
rect 20916 5414 22816 5466
rect 1104 5392 22816 5414
rect 18230 5284 18236 5296
rect 16776 5256 18236 5284
rect 16776 5225 16804 5256
rect 18230 5244 18236 5256
rect 18288 5244 18294 5296
rect 16761 5219 16819 5225
rect 16761 5185 16773 5219
rect 16807 5185 16819 5219
rect 16761 5179 16819 5185
rect 16850 5176 16856 5228
rect 16908 5176 16914 5228
rect 16942 5108 16948 5160
rect 17000 5108 17006 5160
rect 17126 4972 17132 5024
rect 17184 4972 17190 5024
rect 1104 4922 22816 4944
rect 1104 4870 3664 4922
rect 3716 4870 3728 4922
rect 3780 4870 3792 4922
rect 3844 4870 3856 4922
rect 3908 4870 3920 4922
rect 3972 4870 9092 4922
rect 9144 4870 9156 4922
rect 9208 4870 9220 4922
rect 9272 4870 9284 4922
rect 9336 4870 9348 4922
rect 9400 4870 14520 4922
rect 14572 4870 14584 4922
rect 14636 4870 14648 4922
rect 14700 4870 14712 4922
rect 14764 4870 14776 4922
rect 14828 4870 19948 4922
rect 20000 4870 20012 4922
rect 20064 4870 20076 4922
rect 20128 4870 20140 4922
rect 20192 4870 20204 4922
rect 20256 4870 22816 4922
rect 1104 4848 22816 4870
rect 1104 4378 22816 4400
rect 1104 4326 4324 4378
rect 4376 4326 4388 4378
rect 4440 4326 4452 4378
rect 4504 4326 4516 4378
rect 4568 4326 4580 4378
rect 4632 4326 9752 4378
rect 9804 4326 9816 4378
rect 9868 4326 9880 4378
rect 9932 4326 9944 4378
rect 9996 4326 10008 4378
rect 10060 4326 15180 4378
rect 15232 4326 15244 4378
rect 15296 4326 15308 4378
rect 15360 4326 15372 4378
rect 15424 4326 15436 4378
rect 15488 4326 20608 4378
rect 20660 4326 20672 4378
rect 20724 4326 20736 4378
rect 20788 4326 20800 4378
rect 20852 4326 20864 4378
rect 20916 4326 22816 4378
rect 1104 4304 22816 4326
rect 4632 4168 4844 4196
rect 4062 4088 4068 4140
rect 4120 4128 4126 4140
rect 4632 4128 4660 4168
rect 4120 4100 4660 4128
rect 4120 4088 4126 4100
rect 4706 4088 4712 4140
rect 4764 4088 4770 4140
rect 4816 4128 4844 4168
rect 7944 4168 8340 4196
rect 7944 4128 7972 4168
rect 4816 4100 7972 4128
rect 8018 4088 8024 4140
rect 8076 4128 8082 4140
rect 8202 4128 8208 4140
rect 8076 4100 8208 4128
rect 8076 4088 8082 4100
rect 8202 4088 8208 4100
rect 8260 4088 8266 4140
rect 8312 4137 8340 4168
rect 18138 4156 18144 4208
rect 18196 4156 18202 4208
rect 8297 4131 8355 4137
rect 8297 4097 8309 4131
rect 8343 4097 8355 4131
rect 8297 4091 8355 4097
rect 8386 4088 8392 4140
rect 8444 4128 8450 4140
rect 16942 4128 16948 4140
rect 8444 4100 16948 4128
rect 8444 4088 8450 4100
rect 16942 4088 16948 4100
rect 17000 4128 17006 4140
rect 18156 4128 18184 4156
rect 22094 4128 22100 4140
rect 17000 4100 22100 4128
rect 17000 4088 17006 4100
rect 22094 4088 22100 4100
rect 22152 4088 22158 4140
rect 4724 4060 4752 4088
rect 8113 4063 8171 4069
rect 8113 4060 8125 4063
rect 4724 4032 8125 4060
rect 8113 4029 8125 4032
rect 8159 4060 8171 4063
rect 16850 4060 16856 4072
rect 8159 4032 8248 4060
rect 8159 4029 8171 4032
rect 8113 4023 8171 4029
rect 8220 3992 8248 4032
rect 12406 4032 16856 4060
rect 12406 3992 12434 4032
rect 16850 4020 16856 4032
rect 16908 4020 16914 4072
rect 8220 3964 12434 3992
rect 8478 3884 8484 3936
rect 8536 3884 8542 3936
rect 1104 3834 22816 3856
rect 1104 3782 3664 3834
rect 3716 3782 3728 3834
rect 3780 3782 3792 3834
rect 3844 3782 3856 3834
rect 3908 3782 3920 3834
rect 3972 3782 9092 3834
rect 9144 3782 9156 3834
rect 9208 3782 9220 3834
rect 9272 3782 9284 3834
rect 9336 3782 9348 3834
rect 9400 3782 14520 3834
rect 14572 3782 14584 3834
rect 14636 3782 14648 3834
rect 14700 3782 14712 3834
rect 14764 3782 14776 3834
rect 14828 3782 19948 3834
rect 20000 3782 20012 3834
rect 20064 3782 20076 3834
rect 20128 3782 20140 3834
rect 20192 3782 20204 3834
rect 20256 3782 22816 3834
rect 1104 3760 22816 3782
rect 1104 3290 22816 3312
rect 1104 3238 4324 3290
rect 4376 3238 4388 3290
rect 4440 3238 4452 3290
rect 4504 3238 4516 3290
rect 4568 3238 4580 3290
rect 4632 3238 9752 3290
rect 9804 3238 9816 3290
rect 9868 3238 9880 3290
rect 9932 3238 9944 3290
rect 9996 3238 10008 3290
rect 10060 3238 15180 3290
rect 15232 3238 15244 3290
rect 15296 3238 15308 3290
rect 15360 3238 15372 3290
rect 15424 3238 15436 3290
rect 15488 3238 20608 3290
rect 20660 3238 20672 3290
rect 20724 3238 20736 3290
rect 20788 3238 20800 3290
rect 20852 3238 20864 3290
rect 20916 3238 22816 3290
rect 1104 3216 22816 3238
rect 1104 2746 22816 2768
rect 1104 2694 3664 2746
rect 3716 2694 3728 2746
rect 3780 2694 3792 2746
rect 3844 2694 3856 2746
rect 3908 2694 3920 2746
rect 3972 2694 9092 2746
rect 9144 2694 9156 2746
rect 9208 2694 9220 2746
rect 9272 2694 9284 2746
rect 9336 2694 9348 2746
rect 9400 2694 14520 2746
rect 14572 2694 14584 2746
rect 14636 2694 14648 2746
rect 14700 2694 14712 2746
rect 14764 2694 14776 2746
rect 14828 2694 19948 2746
rect 20000 2694 20012 2746
rect 20064 2694 20076 2746
rect 20128 2694 20140 2746
rect 20192 2694 20204 2746
rect 20256 2694 22816 2746
rect 1104 2672 22816 2694
rect 1765 2635 1823 2641
rect 1765 2601 1777 2635
rect 1811 2632 1823 2635
rect 4706 2632 4712 2644
rect 1811 2604 4712 2632
rect 1811 2601 1823 2604
rect 1765 2595 1823 2601
rect 4706 2592 4712 2604
rect 4764 2592 4770 2644
rect 22094 2592 22100 2644
rect 22152 2592 22158 2644
rect 8478 2388 8484 2440
rect 8536 2428 8542 2440
rect 9033 2431 9091 2437
rect 9033 2428 9045 2431
rect 8536 2400 9045 2428
rect 8536 2388 8542 2400
rect 9033 2397 9045 2400
rect 9079 2397 9091 2431
rect 9033 2391 9091 2397
rect 16945 2431 17003 2437
rect 16945 2397 16957 2431
rect 16991 2428 17003 2431
rect 17126 2428 17132 2440
rect 16991 2400 17132 2428
rect 16991 2397 17003 2400
rect 16945 2391 17003 2397
rect 17126 2388 17132 2400
rect 17184 2388 17190 2440
rect 14 2320 20 2372
rect 72 2360 78 2372
rect 1489 2363 1547 2369
rect 1489 2360 1501 2363
rect 72 2332 1501 2360
rect 72 2320 78 2332
rect 1489 2329 1501 2332
rect 1535 2329 1547 2363
rect 1489 2323 1547 2329
rect 22373 2363 22431 2369
rect 22373 2329 22385 2363
rect 22419 2360 22431 2363
rect 22830 2360 22836 2372
rect 22419 2332 22836 2360
rect 22419 2329 22431 2332
rect 22373 2323 22431 2329
rect 22830 2320 22836 2332
rect 22888 2320 22894 2372
rect 8386 2252 8392 2304
rect 8444 2292 8450 2304
rect 9125 2295 9183 2301
rect 9125 2292 9137 2295
rect 8444 2264 9137 2292
rect 8444 2252 8450 2264
rect 9125 2261 9137 2264
rect 9171 2261 9183 2295
rect 9125 2255 9183 2261
rect 16758 2252 16764 2304
rect 16816 2292 16822 2304
rect 17037 2295 17095 2301
rect 17037 2292 17049 2295
rect 16816 2264 17049 2292
rect 16816 2252 16822 2264
rect 17037 2261 17049 2264
rect 17083 2261 17095 2295
rect 17037 2255 17095 2261
rect 1104 2202 22816 2224
rect 1104 2150 4324 2202
rect 4376 2150 4388 2202
rect 4440 2150 4452 2202
rect 4504 2150 4516 2202
rect 4568 2150 4580 2202
rect 4632 2150 9752 2202
rect 9804 2150 9816 2202
rect 9868 2150 9880 2202
rect 9932 2150 9944 2202
rect 9996 2150 10008 2202
rect 10060 2150 15180 2202
rect 15232 2150 15244 2202
rect 15296 2150 15308 2202
rect 15360 2150 15372 2202
rect 15424 2150 15436 2202
rect 15488 2150 20608 2202
rect 20660 2150 20672 2202
rect 20724 2150 20736 2202
rect 20788 2150 20800 2202
rect 20852 2150 20864 2202
rect 20916 2150 22816 2202
rect 1104 2128 22816 2150
<< via1 >>
rect 4324 21734 4376 21786
rect 4388 21734 4440 21786
rect 4452 21734 4504 21786
rect 4516 21734 4568 21786
rect 4580 21734 4632 21786
rect 9752 21734 9804 21786
rect 9816 21734 9868 21786
rect 9880 21734 9932 21786
rect 9944 21734 9996 21786
rect 10008 21734 10060 21786
rect 15180 21734 15232 21786
rect 15244 21734 15296 21786
rect 15308 21734 15360 21786
rect 15372 21734 15424 21786
rect 15436 21734 15488 21786
rect 20608 21734 20660 21786
rect 20672 21734 20724 21786
rect 20736 21734 20788 21786
rect 20800 21734 20852 21786
rect 20864 21734 20916 21786
rect 2596 21675 2648 21684
rect 2596 21641 2605 21675
rect 2605 21641 2639 21675
rect 2639 21641 2648 21675
rect 2596 21632 2648 21641
rect 11152 21632 11204 21684
rect 20260 21675 20312 21684
rect 20260 21641 20269 21675
rect 20269 21641 20303 21675
rect 20303 21641 20312 21675
rect 20260 21632 20312 21641
rect 4252 21496 4304 21548
rect 10968 21496 11020 21548
rect 18052 21496 18104 21548
rect 3664 21190 3716 21242
rect 3728 21190 3780 21242
rect 3792 21190 3844 21242
rect 3856 21190 3908 21242
rect 3920 21190 3972 21242
rect 9092 21190 9144 21242
rect 9156 21190 9208 21242
rect 9220 21190 9272 21242
rect 9284 21190 9336 21242
rect 9348 21190 9400 21242
rect 14520 21190 14572 21242
rect 14584 21190 14636 21242
rect 14648 21190 14700 21242
rect 14712 21190 14764 21242
rect 14776 21190 14828 21242
rect 19948 21190 20000 21242
rect 20012 21190 20064 21242
rect 20076 21190 20128 21242
rect 20140 21190 20192 21242
rect 20204 21190 20256 21242
rect 4324 20646 4376 20698
rect 4388 20646 4440 20698
rect 4452 20646 4504 20698
rect 4516 20646 4568 20698
rect 4580 20646 4632 20698
rect 9752 20646 9804 20698
rect 9816 20646 9868 20698
rect 9880 20646 9932 20698
rect 9944 20646 9996 20698
rect 10008 20646 10060 20698
rect 15180 20646 15232 20698
rect 15244 20646 15296 20698
rect 15308 20646 15360 20698
rect 15372 20646 15424 20698
rect 15436 20646 15488 20698
rect 20608 20646 20660 20698
rect 20672 20646 20724 20698
rect 20736 20646 20788 20698
rect 20800 20646 20852 20698
rect 20864 20646 20916 20698
rect 3664 20102 3716 20154
rect 3728 20102 3780 20154
rect 3792 20102 3844 20154
rect 3856 20102 3908 20154
rect 3920 20102 3972 20154
rect 9092 20102 9144 20154
rect 9156 20102 9208 20154
rect 9220 20102 9272 20154
rect 9284 20102 9336 20154
rect 9348 20102 9400 20154
rect 14520 20102 14572 20154
rect 14584 20102 14636 20154
rect 14648 20102 14700 20154
rect 14712 20102 14764 20154
rect 14776 20102 14828 20154
rect 19948 20102 20000 20154
rect 20012 20102 20064 20154
rect 20076 20102 20128 20154
rect 20140 20102 20192 20154
rect 20204 20102 20256 20154
rect 22836 19932 22888 19984
rect 22192 19839 22244 19848
rect 22192 19805 22201 19839
rect 22201 19805 22235 19839
rect 22235 19805 22244 19839
rect 22192 19796 22244 19805
rect 4324 19558 4376 19610
rect 4388 19558 4440 19610
rect 4452 19558 4504 19610
rect 4516 19558 4568 19610
rect 4580 19558 4632 19610
rect 9752 19558 9804 19610
rect 9816 19558 9868 19610
rect 9880 19558 9932 19610
rect 9944 19558 9996 19610
rect 10008 19558 10060 19610
rect 15180 19558 15232 19610
rect 15244 19558 15296 19610
rect 15308 19558 15360 19610
rect 15372 19558 15424 19610
rect 15436 19558 15488 19610
rect 20608 19558 20660 19610
rect 20672 19558 20724 19610
rect 20736 19558 20788 19610
rect 20800 19558 20852 19610
rect 20864 19558 20916 19610
rect 3664 19014 3716 19066
rect 3728 19014 3780 19066
rect 3792 19014 3844 19066
rect 3856 19014 3908 19066
rect 3920 19014 3972 19066
rect 9092 19014 9144 19066
rect 9156 19014 9208 19066
rect 9220 19014 9272 19066
rect 9284 19014 9336 19066
rect 9348 19014 9400 19066
rect 14520 19014 14572 19066
rect 14584 19014 14636 19066
rect 14648 19014 14700 19066
rect 14712 19014 14764 19066
rect 14776 19014 14828 19066
rect 19948 19014 20000 19066
rect 20012 19014 20064 19066
rect 20076 19014 20128 19066
rect 20140 19014 20192 19066
rect 20204 19014 20256 19066
rect 4252 18955 4304 18964
rect 4252 18921 4261 18955
rect 4261 18921 4295 18955
rect 4295 18921 4304 18955
rect 4252 18912 4304 18921
rect 10968 18955 11020 18964
rect 10968 18921 10977 18955
rect 10977 18921 11011 18955
rect 11011 18921 11020 18955
rect 10968 18912 11020 18921
rect 4252 18708 4304 18760
rect 10784 18751 10836 18760
rect 10784 18717 10793 18751
rect 10793 18717 10827 18751
rect 10827 18717 10836 18751
rect 10784 18708 10836 18717
rect 4324 18470 4376 18522
rect 4388 18470 4440 18522
rect 4452 18470 4504 18522
rect 4516 18470 4568 18522
rect 4580 18470 4632 18522
rect 9752 18470 9804 18522
rect 9816 18470 9868 18522
rect 9880 18470 9932 18522
rect 9944 18470 9996 18522
rect 10008 18470 10060 18522
rect 15180 18470 15232 18522
rect 15244 18470 15296 18522
rect 15308 18470 15360 18522
rect 15372 18470 15424 18522
rect 15436 18470 15488 18522
rect 20608 18470 20660 18522
rect 20672 18470 20724 18522
rect 20736 18470 20788 18522
rect 20800 18470 20852 18522
rect 20864 18470 20916 18522
rect 4252 18411 4304 18420
rect 4252 18377 4261 18411
rect 4261 18377 4295 18411
rect 4295 18377 4304 18411
rect 4252 18368 4304 18377
rect 10784 18368 10836 18420
rect 22192 18368 22244 18420
rect 4160 18300 4212 18352
rect 1492 18275 1544 18284
rect 1492 18241 1501 18275
rect 1501 18241 1535 18275
rect 1535 18241 1544 18275
rect 1492 18232 1544 18241
rect 18972 18275 19024 18284
rect 18972 18241 18981 18275
rect 18981 18241 19015 18275
rect 19015 18241 19024 18275
rect 18972 18232 19024 18241
rect 4068 18028 4120 18080
rect 15200 18096 15252 18148
rect 17500 18028 17552 18080
rect 3664 17926 3716 17978
rect 3728 17926 3780 17978
rect 3792 17926 3844 17978
rect 3856 17926 3908 17978
rect 3920 17926 3972 17978
rect 9092 17926 9144 17978
rect 9156 17926 9208 17978
rect 9220 17926 9272 17978
rect 9284 17926 9336 17978
rect 9348 17926 9400 17978
rect 14520 17926 14572 17978
rect 14584 17926 14636 17978
rect 14648 17926 14700 17978
rect 14712 17926 14764 17978
rect 14776 17926 14828 17978
rect 19948 17926 20000 17978
rect 20012 17926 20064 17978
rect 20076 17926 20128 17978
rect 20140 17926 20192 17978
rect 20204 17926 20256 17978
rect 18052 17824 18104 17876
rect 18144 17867 18196 17876
rect 18144 17833 18153 17867
rect 18153 17833 18187 17867
rect 18187 17833 18196 17867
rect 18144 17824 18196 17833
rect 18972 17824 19024 17876
rect 17500 17799 17552 17808
rect 17500 17765 17509 17799
rect 17509 17765 17543 17799
rect 17543 17765 17552 17799
rect 17500 17756 17552 17765
rect 15200 17688 15252 17740
rect 17776 17663 17828 17672
rect 17776 17629 17785 17663
rect 17785 17629 17819 17663
rect 17819 17629 17828 17663
rect 17776 17620 17828 17629
rect 18236 17484 18288 17536
rect 4324 17382 4376 17434
rect 4388 17382 4440 17434
rect 4452 17382 4504 17434
rect 4516 17382 4568 17434
rect 4580 17382 4632 17434
rect 9752 17382 9804 17434
rect 9816 17382 9868 17434
rect 9880 17382 9932 17434
rect 9944 17382 9996 17434
rect 10008 17382 10060 17434
rect 15180 17382 15232 17434
rect 15244 17382 15296 17434
rect 15308 17382 15360 17434
rect 15372 17382 15424 17434
rect 15436 17382 15488 17434
rect 20608 17382 20660 17434
rect 20672 17382 20724 17434
rect 20736 17382 20788 17434
rect 20800 17382 20852 17434
rect 20864 17382 20916 17434
rect 3664 16838 3716 16890
rect 3728 16838 3780 16890
rect 3792 16838 3844 16890
rect 3856 16838 3908 16890
rect 3920 16838 3972 16890
rect 9092 16838 9144 16890
rect 9156 16838 9208 16890
rect 9220 16838 9272 16890
rect 9284 16838 9336 16890
rect 9348 16838 9400 16890
rect 14520 16838 14572 16890
rect 14584 16838 14636 16890
rect 14648 16838 14700 16890
rect 14712 16838 14764 16890
rect 14776 16838 14828 16890
rect 19948 16838 20000 16890
rect 20012 16838 20064 16890
rect 20076 16838 20128 16890
rect 20140 16838 20192 16890
rect 20204 16838 20256 16890
rect 4324 16294 4376 16346
rect 4388 16294 4440 16346
rect 4452 16294 4504 16346
rect 4516 16294 4568 16346
rect 4580 16294 4632 16346
rect 9752 16294 9804 16346
rect 9816 16294 9868 16346
rect 9880 16294 9932 16346
rect 9944 16294 9996 16346
rect 10008 16294 10060 16346
rect 15180 16294 15232 16346
rect 15244 16294 15296 16346
rect 15308 16294 15360 16346
rect 15372 16294 15424 16346
rect 15436 16294 15488 16346
rect 20608 16294 20660 16346
rect 20672 16294 20724 16346
rect 20736 16294 20788 16346
rect 20800 16294 20852 16346
rect 20864 16294 20916 16346
rect 3664 15750 3716 15802
rect 3728 15750 3780 15802
rect 3792 15750 3844 15802
rect 3856 15750 3908 15802
rect 3920 15750 3972 15802
rect 9092 15750 9144 15802
rect 9156 15750 9208 15802
rect 9220 15750 9272 15802
rect 9284 15750 9336 15802
rect 9348 15750 9400 15802
rect 14520 15750 14572 15802
rect 14584 15750 14636 15802
rect 14648 15750 14700 15802
rect 14712 15750 14764 15802
rect 14776 15750 14828 15802
rect 19948 15750 20000 15802
rect 20012 15750 20064 15802
rect 20076 15750 20128 15802
rect 20140 15750 20192 15802
rect 20204 15750 20256 15802
rect 4324 15206 4376 15258
rect 4388 15206 4440 15258
rect 4452 15206 4504 15258
rect 4516 15206 4568 15258
rect 4580 15206 4632 15258
rect 9752 15206 9804 15258
rect 9816 15206 9868 15258
rect 9880 15206 9932 15258
rect 9944 15206 9996 15258
rect 10008 15206 10060 15258
rect 15180 15206 15232 15258
rect 15244 15206 15296 15258
rect 15308 15206 15360 15258
rect 15372 15206 15424 15258
rect 15436 15206 15488 15258
rect 20608 15206 20660 15258
rect 20672 15206 20724 15258
rect 20736 15206 20788 15258
rect 20800 15206 20852 15258
rect 20864 15206 20916 15258
rect 3664 14662 3716 14714
rect 3728 14662 3780 14714
rect 3792 14662 3844 14714
rect 3856 14662 3908 14714
rect 3920 14662 3972 14714
rect 9092 14662 9144 14714
rect 9156 14662 9208 14714
rect 9220 14662 9272 14714
rect 9284 14662 9336 14714
rect 9348 14662 9400 14714
rect 14520 14662 14572 14714
rect 14584 14662 14636 14714
rect 14648 14662 14700 14714
rect 14712 14662 14764 14714
rect 14776 14662 14828 14714
rect 19948 14662 20000 14714
rect 20012 14662 20064 14714
rect 20076 14662 20128 14714
rect 20140 14662 20192 14714
rect 20204 14662 20256 14714
rect 4324 14118 4376 14170
rect 4388 14118 4440 14170
rect 4452 14118 4504 14170
rect 4516 14118 4568 14170
rect 4580 14118 4632 14170
rect 9752 14118 9804 14170
rect 9816 14118 9868 14170
rect 9880 14118 9932 14170
rect 9944 14118 9996 14170
rect 10008 14118 10060 14170
rect 15180 14118 15232 14170
rect 15244 14118 15296 14170
rect 15308 14118 15360 14170
rect 15372 14118 15424 14170
rect 15436 14118 15488 14170
rect 20608 14118 20660 14170
rect 20672 14118 20724 14170
rect 20736 14118 20788 14170
rect 20800 14118 20852 14170
rect 20864 14118 20916 14170
rect 3664 13574 3716 13626
rect 3728 13574 3780 13626
rect 3792 13574 3844 13626
rect 3856 13574 3908 13626
rect 3920 13574 3972 13626
rect 9092 13574 9144 13626
rect 9156 13574 9208 13626
rect 9220 13574 9272 13626
rect 9284 13574 9336 13626
rect 9348 13574 9400 13626
rect 14520 13574 14572 13626
rect 14584 13574 14636 13626
rect 14648 13574 14700 13626
rect 14712 13574 14764 13626
rect 14776 13574 14828 13626
rect 19948 13574 20000 13626
rect 20012 13574 20064 13626
rect 20076 13574 20128 13626
rect 20140 13574 20192 13626
rect 20204 13574 20256 13626
rect 4324 13030 4376 13082
rect 4388 13030 4440 13082
rect 4452 13030 4504 13082
rect 4516 13030 4568 13082
rect 4580 13030 4632 13082
rect 9752 13030 9804 13082
rect 9816 13030 9868 13082
rect 9880 13030 9932 13082
rect 9944 13030 9996 13082
rect 10008 13030 10060 13082
rect 15180 13030 15232 13082
rect 15244 13030 15296 13082
rect 15308 13030 15360 13082
rect 15372 13030 15424 13082
rect 15436 13030 15488 13082
rect 20608 13030 20660 13082
rect 20672 13030 20724 13082
rect 20736 13030 20788 13082
rect 20800 13030 20852 13082
rect 20864 13030 20916 13082
rect 3664 12486 3716 12538
rect 3728 12486 3780 12538
rect 3792 12486 3844 12538
rect 3856 12486 3908 12538
rect 3920 12486 3972 12538
rect 9092 12486 9144 12538
rect 9156 12486 9208 12538
rect 9220 12486 9272 12538
rect 9284 12486 9336 12538
rect 9348 12486 9400 12538
rect 14520 12486 14572 12538
rect 14584 12486 14636 12538
rect 14648 12486 14700 12538
rect 14712 12486 14764 12538
rect 14776 12486 14828 12538
rect 19948 12486 20000 12538
rect 20012 12486 20064 12538
rect 20076 12486 20128 12538
rect 20140 12486 20192 12538
rect 20204 12486 20256 12538
rect 4324 11942 4376 11994
rect 4388 11942 4440 11994
rect 4452 11942 4504 11994
rect 4516 11942 4568 11994
rect 4580 11942 4632 11994
rect 9752 11942 9804 11994
rect 9816 11942 9868 11994
rect 9880 11942 9932 11994
rect 9944 11942 9996 11994
rect 10008 11942 10060 11994
rect 15180 11942 15232 11994
rect 15244 11942 15296 11994
rect 15308 11942 15360 11994
rect 15372 11942 15424 11994
rect 15436 11942 15488 11994
rect 20608 11942 20660 11994
rect 20672 11942 20724 11994
rect 20736 11942 20788 11994
rect 20800 11942 20852 11994
rect 20864 11942 20916 11994
rect 3664 11398 3716 11450
rect 3728 11398 3780 11450
rect 3792 11398 3844 11450
rect 3856 11398 3908 11450
rect 3920 11398 3972 11450
rect 9092 11398 9144 11450
rect 9156 11398 9208 11450
rect 9220 11398 9272 11450
rect 9284 11398 9336 11450
rect 9348 11398 9400 11450
rect 14520 11398 14572 11450
rect 14584 11398 14636 11450
rect 14648 11398 14700 11450
rect 14712 11398 14764 11450
rect 14776 11398 14828 11450
rect 19948 11398 20000 11450
rect 20012 11398 20064 11450
rect 20076 11398 20128 11450
rect 20140 11398 20192 11450
rect 20204 11398 20256 11450
rect 4324 10854 4376 10906
rect 4388 10854 4440 10906
rect 4452 10854 4504 10906
rect 4516 10854 4568 10906
rect 4580 10854 4632 10906
rect 9752 10854 9804 10906
rect 9816 10854 9868 10906
rect 9880 10854 9932 10906
rect 9944 10854 9996 10906
rect 10008 10854 10060 10906
rect 15180 10854 15232 10906
rect 15244 10854 15296 10906
rect 15308 10854 15360 10906
rect 15372 10854 15424 10906
rect 15436 10854 15488 10906
rect 20608 10854 20660 10906
rect 20672 10854 20724 10906
rect 20736 10854 20788 10906
rect 20800 10854 20852 10906
rect 20864 10854 20916 10906
rect 18880 10659 18932 10668
rect 18880 10625 18889 10659
rect 18889 10625 18923 10659
rect 18923 10625 18932 10659
rect 18880 10616 18932 10625
rect 22376 10455 22428 10464
rect 22376 10421 22385 10455
rect 22385 10421 22419 10455
rect 22419 10421 22428 10455
rect 22376 10412 22428 10421
rect 3664 10310 3716 10362
rect 3728 10310 3780 10362
rect 3792 10310 3844 10362
rect 3856 10310 3908 10362
rect 3920 10310 3972 10362
rect 9092 10310 9144 10362
rect 9156 10310 9208 10362
rect 9220 10310 9272 10362
rect 9284 10310 9336 10362
rect 9348 10310 9400 10362
rect 14520 10310 14572 10362
rect 14584 10310 14636 10362
rect 14648 10310 14700 10362
rect 14712 10310 14764 10362
rect 14776 10310 14828 10362
rect 19948 10310 20000 10362
rect 20012 10310 20064 10362
rect 20076 10310 20128 10362
rect 20140 10310 20192 10362
rect 20204 10310 20256 10362
rect 18144 10251 18196 10260
rect 18144 10217 18153 10251
rect 18153 10217 18187 10251
rect 18187 10217 18196 10251
rect 18144 10208 18196 10217
rect 18880 10208 18932 10260
rect 18236 10004 18288 10056
rect 16856 9936 16908 9988
rect 17776 9936 17828 9988
rect 4324 9766 4376 9818
rect 4388 9766 4440 9818
rect 4452 9766 4504 9818
rect 4516 9766 4568 9818
rect 4580 9766 4632 9818
rect 9752 9766 9804 9818
rect 9816 9766 9868 9818
rect 9880 9766 9932 9818
rect 9944 9766 9996 9818
rect 10008 9766 10060 9818
rect 15180 9766 15232 9818
rect 15244 9766 15296 9818
rect 15308 9766 15360 9818
rect 15372 9766 15424 9818
rect 15436 9766 15488 9818
rect 20608 9766 20660 9818
rect 20672 9766 20724 9818
rect 20736 9766 20788 9818
rect 20800 9766 20852 9818
rect 20864 9766 20916 9818
rect 3664 9222 3716 9274
rect 3728 9222 3780 9274
rect 3792 9222 3844 9274
rect 3856 9222 3908 9274
rect 3920 9222 3972 9274
rect 9092 9222 9144 9274
rect 9156 9222 9208 9274
rect 9220 9222 9272 9274
rect 9284 9222 9336 9274
rect 9348 9222 9400 9274
rect 14520 9222 14572 9274
rect 14584 9222 14636 9274
rect 14648 9222 14700 9274
rect 14712 9222 14764 9274
rect 14776 9222 14828 9274
rect 19948 9222 20000 9274
rect 20012 9222 20064 9274
rect 20076 9222 20128 9274
rect 20140 9222 20192 9274
rect 20204 9222 20256 9274
rect 4160 9027 4212 9036
rect 4160 8993 4169 9027
rect 4169 8993 4203 9027
rect 4203 8993 4212 9027
rect 4160 8984 4212 8993
rect 4712 8984 4764 9036
rect 4068 8959 4120 8968
rect 4068 8925 4077 8959
rect 4077 8925 4111 8959
rect 4111 8925 4120 8959
rect 4068 8916 4120 8925
rect 8024 8916 8076 8968
rect 940 8848 992 8900
rect 4324 8678 4376 8730
rect 4388 8678 4440 8730
rect 4452 8678 4504 8730
rect 4516 8678 4568 8730
rect 4580 8678 4632 8730
rect 9752 8678 9804 8730
rect 9816 8678 9868 8730
rect 9880 8678 9932 8730
rect 9944 8678 9996 8730
rect 10008 8678 10060 8730
rect 15180 8678 15232 8730
rect 15244 8678 15296 8730
rect 15308 8678 15360 8730
rect 15372 8678 15424 8730
rect 15436 8678 15488 8730
rect 20608 8678 20660 8730
rect 20672 8678 20724 8730
rect 20736 8678 20788 8730
rect 20800 8678 20852 8730
rect 20864 8678 20916 8730
rect 3664 8134 3716 8186
rect 3728 8134 3780 8186
rect 3792 8134 3844 8186
rect 3856 8134 3908 8186
rect 3920 8134 3972 8186
rect 9092 8134 9144 8186
rect 9156 8134 9208 8186
rect 9220 8134 9272 8186
rect 9284 8134 9336 8186
rect 9348 8134 9400 8186
rect 14520 8134 14572 8186
rect 14584 8134 14636 8186
rect 14648 8134 14700 8186
rect 14712 8134 14764 8186
rect 14776 8134 14828 8186
rect 19948 8134 20000 8186
rect 20012 8134 20064 8186
rect 20076 8134 20128 8186
rect 20140 8134 20192 8186
rect 20204 8134 20256 8186
rect 4324 7590 4376 7642
rect 4388 7590 4440 7642
rect 4452 7590 4504 7642
rect 4516 7590 4568 7642
rect 4580 7590 4632 7642
rect 9752 7590 9804 7642
rect 9816 7590 9868 7642
rect 9880 7590 9932 7642
rect 9944 7590 9996 7642
rect 10008 7590 10060 7642
rect 15180 7590 15232 7642
rect 15244 7590 15296 7642
rect 15308 7590 15360 7642
rect 15372 7590 15424 7642
rect 15436 7590 15488 7642
rect 20608 7590 20660 7642
rect 20672 7590 20724 7642
rect 20736 7590 20788 7642
rect 20800 7590 20852 7642
rect 20864 7590 20916 7642
rect 3664 7046 3716 7098
rect 3728 7046 3780 7098
rect 3792 7046 3844 7098
rect 3856 7046 3908 7098
rect 3920 7046 3972 7098
rect 9092 7046 9144 7098
rect 9156 7046 9208 7098
rect 9220 7046 9272 7098
rect 9284 7046 9336 7098
rect 9348 7046 9400 7098
rect 14520 7046 14572 7098
rect 14584 7046 14636 7098
rect 14648 7046 14700 7098
rect 14712 7046 14764 7098
rect 14776 7046 14828 7098
rect 19948 7046 20000 7098
rect 20012 7046 20064 7098
rect 20076 7046 20128 7098
rect 20140 7046 20192 7098
rect 20204 7046 20256 7098
rect 4324 6502 4376 6554
rect 4388 6502 4440 6554
rect 4452 6502 4504 6554
rect 4516 6502 4568 6554
rect 4580 6502 4632 6554
rect 9752 6502 9804 6554
rect 9816 6502 9868 6554
rect 9880 6502 9932 6554
rect 9944 6502 9996 6554
rect 10008 6502 10060 6554
rect 15180 6502 15232 6554
rect 15244 6502 15296 6554
rect 15308 6502 15360 6554
rect 15372 6502 15424 6554
rect 15436 6502 15488 6554
rect 20608 6502 20660 6554
rect 20672 6502 20724 6554
rect 20736 6502 20788 6554
rect 20800 6502 20852 6554
rect 20864 6502 20916 6554
rect 3664 5958 3716 6010
rect 3728 5958 3780 6010
rect 3792 5958 3844 6010
rect 3856 5958 3908 6010
rect 3920 5958 3972 6010
rect 9092 5958 9144 6010
rect 9156 5958 9208 6010
rect 9220 5958 9272 6010
rect 9284 5958 9336 6010
rect 9348 5958 9400 6010
rect 14520 5958 14572 6010
rect 14584 5958 14636 6010
rect 14648 5958 14700 6010
rect 14712 5958 14764 6010
rect 14776 5958 14828 6010
rect 19948 5958 20000 6010
rect 20012 5958 20064 6010
rect 20076 5958 20128 6010
rect 20140 5958 20192 6010
rect 20204 5958 20256 6010
rect 4324 5414 4376 5466
rect 4388 5414 4440 5466
rect 4452 5414 4504 5466
rect 4516 5414 4568 5466
rect 4580 5414 4632 5466
rect 9752 5414 9804 5466
rect 9816 5414 9868 5466
rect 9880 5414 9932 5466
rect 9944 5414 9996 5466
rect 10008 5414 10060 5466
rect 15180 5414 15232 5466
rect 15244 5414 15296 5466
rect 15308 5414 15360 5466
rect 15372 5414 15424 5466
rect 15436 5414 15488 5466
rect 20608 5414 20660 5466
rect 20672 5414 20724 5466
rect 20736 5414 20788 5466
rect 20800 5414 20852 5466
rect 20864 5414 20916 5466
rect 18236 5244 18288 5296
rect 16856 5219 16908 5228
rect 16856 5185 16865 5219
rect 16865 5185 16899 5219
rect 16899 5185 16908 5219
rect 16856 5176 16908 5185
rect 16948 5151 17000 5160
rect 16948 5117 16957 5151
rect 16957 5117 16991 5151
rect 16991 5117 17000 5151
rect 16948 5108 17000 5117
rect 17132 5015 17184 5024
rect 17132 4981 17141 5015
rect 17141 4981 17175 5015
rect 17175 4981 17184 5015
rect 17132 4972 17184 4981
rect 3664 4870 3716 4922
rect 3728 4870 3780 4922
rect 3792 4870 3844 4922
rect 3856 4870 3908 4922
rect 3920 4870 3972 4922
rect 9092 4870 9144 4922
rect 9156 4870 9208 4922
rect 9220 4870 9272 4922
rect 9284 4870 9336 4922
rect 9348 4870 9400 4922
rect 14520 4870 14572 4922
rect 14584 4870 14636 4922
rect 14648 4870 14700 4922
rect 14712 4870 14764 4922
rect 14776 4870 14828 4922
rect 19948 4870 20000 4922
rect 20012 4870 20064 4922
rect 20076 4870 20128 4922
rect 20140 4870 20192 4922
rect 20204 4870 20256 4922
rect 4324 4326 4376 4378
rect 4388 4326 4440 4378
rect 4452 4326 4504 4378
rect 4516 4326 4568 4378
rect 4580 4326 4632 4378
rect 9752 4326 9804 4378
rect 9816 4326 9868 4378
rect 9880 4326 9932 4378
rect 9944 4326 9996 4378
rect 10008 4326 10060 4378
rect 15180 4326 15232 4378
rect 15244 4326 15296 4378
rect 15308 4326 15360 4378
rect 15372 4326 15424 4378
rect 15436 4326 15488 4378
rect 20608 4326 20660 4378
rect 20672 4326 20724 4378
rect 20736 4326 20788 4378
rect 20800 4326 20852 4378
rect 20864 4326 20916 4378
rect 4068 4088 4120 4140
rect 4712 4088 4764 4140
rect 8024 4088 8076 4140
rect 8208 4131 8260 4140
rect 8208 4097 8217 4131
rect 8217 4097 8251 4131
rect 8251 4097 8260 4131
rect 8208 4088 8260 4097
rect 18144 4156 18196 4208
rect 8392 4088 8444 4140
rect 16948 4088 17000 4140
rect 22100 4088 22152 4140
rect 16856 4020 16908 4072
rect 8484 3927 8536 3936
rect 8484 3893 8493 3927
rect 8493 3893 8527 3927
rect 8527 3893 8536 3927
rect 8484 3884 8536 3893
rect 3664 3782 3716 3834
rect 3728 3782 3780 3834
rect 3792 3782 3844 3834
rect 3856 3782 3908 3834
rect 3920 3782 3972 3834
rect 9092 3782 9144 3834
rect 9156 3782 9208 3834
rect 9220 3782 9272 3834
rect 9284 3782 9336 3834
rect 9348 3782 9400 3834
rect 14520 3782 14572 3834
rect 14584 3782 14636 3834
rect 14648 3782 14700 3834
rect 14712 3782 14764 3834
rect 14776 3782 14828 3834
rect 19948 3782 20000 3834
rect 20012 3782 20064 3834
rect 20076 3782 20128 3834
rect 20140 3782 20192 3834
rect 20204 3782 20256 3834
rect 4324 3238 4376 3290
rect 4388 3238 4440 3290
rect 4452 3238 4504 3290
rect 4516 3238 4568 3290
rect 4580 3238 4632 3290
rect 9752 3238 9804 3290
rect 9816 3238 9868 3290
rect 9880 3238 9932 3290
rect 9944 3238 9996 3290
rect 10008 3238 10060 3290
rect 15180 3238 15232 3290
rect 15244 3238 15296 3290
rect 15308 3238 15360 3290
rect 15372 3238 15424 3290
rect 15436 3238 15488 3290
rect 20608 3238 20660 3290
rect 20672 3238 20724 3290
rect 20736 3238 20788 3290
rect 20800 3238 20852 3290
rect 20864 3238 20916 3290
rect 3664 2694 3716 2746
rect 3728 2694 3780 2746
rect 3792 2694 3844 2746
rect 3856 2694 3908 2746
rect 3920 2694 3972 2746
rect 9092 2694 9144 2746
rect 9156 2694 9208 2746
rect 9220 2694 9272 2746
rect 9284 2694 9336 2746
rect 9348 2694 9400 2746
rect 14520 2694 14572 2746
rect 14584 2694 14636 2746
rect 14648 2694 14700 2746
rect 14712 2694 14764 2746
rect 14776 2694 14828 2746
rect 19948 2694 20000 2746
rect 20012 2694 20064 2746
rect 20076 2694 20128 2746
rect 20140 2694 20192 2746
rect 20204 2694 20256 2746
rect 4712 2592 4764 2644
rect 22100 2635 22152 2644
rect 22100 2601 22109 2635
rect 22109 2601 22143 2635
rect 22143 2601 22152 2635
rect 22100 2592 22152 2601
rect 8484 2388 8536 2440
rect 17132 2388 17184 2440
rect 20 2320 72 2372
rect 22836 2320 22888 2372
rect 8392 2252 8444 2304
rect 16764 2252 16816 2304
rect 4324 2150 4376 2202
rect 4388 2150 4440 2202
rect 4452 2150 4504 2202
rect 4516 2150 4568 2202
rect 4580 2150 4632 2202
rect 9752 2150 9804 2202
rect 9816 2150 9868 2202
rect 9880 2150 9932 2202
rect 9944 2150 9996 2202
rect 10008 2150 10060 2202
rect 15180 2150 15232 2202
rect 15244 2150 15296 2202
rect 15308 2150 15360 2202
rect 15372 2150 15424 2202
rect 15436 2150 15488 2202
rect 20608 2150 20660 2202
rect 20672 2150 20724 2202
rect 20736 2150 20788 2202
rect 20800 2150 20852 2202
rect 20864 2150 20916 2202
<< metal2 >>
rect 2594 23200 2650 24000
rect 10966 23200 11022 24000
rect 19982 23338 20038 24000
rect 19982 23310 20300 23338
rect 19982 23200 20038 23310
rect 2608 21690 2636 23200
rect 10980 22094 11008 23200
rect 10980 22066 11192 22094
rect 4324 21788 4632 21797
rect 4324 21786 4330 21788
rect 4386 21786 4410 21788
rect 4466 21786 4490 21788
rect 4546 21786 4570 21788
rect 4626 21786 4632 21788
rect 4386 21734 4388 21786
rect 4568 21734 4570 21786
rect 4324 21732 4330 21734
rect 4386 21732 4410 21734
rect 4466 21732 4490 21734
rect 4546 21732 4570 21734
rect 4626 21732 4632 21734
rect 4324 21723 4632 21732
rect 9752 21788 10060 21797
rect 9752 21786 9758 21788
rect 9814 21786 9838 21788
rect 9894 21786 9918 21788
rect 9974 21786 9998 21788
rect 10054 21786 10060 21788
rect 9814 21734 9816 21786
rect 9996 21734 9998 21786
rect 9752 21732 9758 21734
rect 9814 21732 9838 21734
rect 9894 21732 9918 21734
rect 9974 21732 9998 21734
rect 10054 21732 10060 21734
rect 9752 21723 10060 21732
rect 11164 21690 11192 22066
rect 15180 21788 15488 21797
rect 15180 21786 15186 21788
rect 15242 21786 15266 21788
rect 15322 21786 15346 21788
rect 15402 21786 15426 21788
rect 15482 21786 15488 21788
rect 15242 21734 15244 21786
rect 15424 21734 15426 21786
rect 15180 21732 15186 21734
rect 15242 21732 15266 21734
rect 15322 21732 15346 21734
rect 15402 21732 15426 21734
rect 15482 21732 15488 21734
rect 15180 21723 15488 21732
rect 20272 21690 20300 23310
rect 20608 21788 20916 21797
rect 20608 21786 20614 21788
rect 20670 21786 20694 21788
rect 20750 21786 20774 21788
rect 20830 21786 20854 21788
rect 20910 21786 20916 21788
rect 20670 21734 20672 21786
rect 20852 21734 20854 21786
rect 20608 21732 20614 21734
rect 20670 21732 20694 21734
rect 20750 21732 20774 21734
rect 20830 21732 20854 21734
rect 20910 21732 20916 21734
rect 20608 21723 20916 21732
rect 2596 21684 2648 21690
rect 2596 21626 2648 21632
rect 11152 21684 11204 21690
rect 11152 21626 11204 21632
rect 20260 21684 20312 21690
rect 20260 21626 20312 21632
rect 4252 21548 4304 21554
rect 4252 21490 4304 21496
rect 10968 21548 11020 21554
rect 10968 21490 11020 21496
rect 18052 21548 18104 21554
rect 18052 21490 18104 21496
rect 3664 21244 3972 21253
rect 3664 21242 3670 21244
rect 3726 21242 3750 21244
rect 3806 21242 3830 21244
rect 3886 21242 3910 21244
rect 3966 21242 3972 21244
rect 3726 21190 3728 21242
rect 3908 21190 3910 21242
rect 3664 21188 3670 21190
rect 3726 21188 3750 21190
rect 3806 21188 3830 21190
rect 3886 21188 3910 21190
rect 3966 21188 3972 21190
rect 3664 21179 3972 21188
rect 3664 20156 3972 20165
rect 3664 20154 3670 20156
rect 3726 20154 3750 20156
rect 3806 20154 3830 20156
rect 3886 20154 3910 20156
rect 3966 20154 3972 20156
rect 3726 20102 3728 20154
rect 3908 20102 3910 20154
rect 3664 20100 3670 20102
rect 3726 20100 3750 20102
rect 3806 20100 3830 20102
rect 3886 20100 3910 20102
rect 3966 20100 3972 20102
rect 3664 20091 3972 20100
rect 3664 19068 3972 19077
rect 3664 19066 3670 19068
rect 3726 19066 3750 19068
rect 3806 19066 3830 19068
rect 3886 19066 3910 19068
rect 3966 19066 3972 19068
rect 3726 19014 3728 19066
rect 3908 19014 3910 19066
rect 3664 19012 3670 19014
rect 3726 19012 3750 19014
rect 3806 19012 3830 19014
rect 3886 19012 3910 19014
rect 3966 19012 3972 19014
rect 3664 19003 3972 19012
rect 4264 18970 4292 21490
rect 9092 21244 9400 21253
rect 9092 21242 9098 21244
rect 9154 21242 9178 21244
rect 9234 21242 9258 21244
rect 9314 21242 9338 21244
rect 9394 21242 9400 21244
rect 9154 21190 9156 21242
rect 9336 21190 9338 21242
rect 9092 21188 9098 21190
rect 9154 21188 9178 21190
rect 9234 21188 9258 21190
rect 9314 21188 9338 21190
rect 9394 21188 9400 21190
rect 9092 21179 9400 21188
rect 4324 20700 4632 20709
rect 4324 20698 4330 20700
rect 4386 20698 4410 20700
rect 4466 20698 4490 20700
rect 4546 20698 4570 20700
rect 4626 20698 4632 20700
rect 4386 20646 4388 20698
rect 4568 20646 4570 20698
rect 4324 20644 4330 20646
rect 4386 20644 4410 20646
rect 4466 20644 4490 20646
rect 4546 20644 4570 20646
rect 4626 20644 4632 20646
rect 4324 20635 4632 20644
rect 9752 20700 10060 20709
rect 9752 20698 9758 20700
rect 9814 20698 9838 20700
rect 9894 20698 9918 20700
rect 9974 20698 9998 20700
rect 10054 20698 10060 20700
rect 9814 20646 9816 20698
rect 9996 20646 9998 20698
rect 9752 20644 9758 20646
rect 9814 20644 9838 20646
rect 9894 20644 9918 20646
rect 9974 20644 9998 20646
rect 10054 20644 10060 20646
rect 9752 20635 10060 20644
rect 9092 20156 9400 20165
rect 9092 20154 9098 20156
rect 9154 20154 9178 20156
rect 9234 20154 9258 20156
rect 9314 20154 9338 20156
rect 9394 20154 9400 20156
rect 9154 20102 9156 20154
rect 9336 20102 9338 20154
rect 9092 20100 9098 20102
rect 9154 20100 9178 20102
rect 9234 20100 9258 20102
rect 9314 20100 9338 20102
rect 9394 20100 9400 20102
rect 9092 20091 9400 20100
rect 4324 19612 4632 19621
rect 4324 19610 4330 19612
rect 4386 19610 4410 19612
rect 4466 19610 4490 19612
rect 4546 19610 4570 19612
rect 4626 19610 4632 19612
rect 4386 19558 4388 19610
rect 4568 19558 4570 19610
rect 4324 19556 4330 19558
rect 4386 19556 4410 19558
rect 4466 19556 4490 19558
rect 4546 19556 4570 19558
rect 4626 19556 4632 19558
rect 4324 19547 4632 19556
rect 9752 19612 10060 19621
rect 9752 19610 9758 19612
rect 9814 19610 9838 19612
rect 9894 19610 9918 19612
rect 9974 19610 9998 19612
rect 10054 19610 10060 19612
rect 9814 19558 9816 19610
rect 9996 19558 9998 19610
rect 9752 19556 9758 19558
rect 9814 19556 9838 19558
rect 9894 19556 9918 19558
rect 9974 19556 9998 19558
rect 10054 19556 10060 19558
rect 9752 19547 10060 19556
rect 9092 19068 9400 19077
rect 9092 19066 9098 19068
rect 9154 19066 9178 19068
rect 9234 19066 9258 19068
rect 9314 19066 9338 19068
rect 9394 19066 9400 19068
rect 9154 19014 9156 19066
rect 9336 19014 9338 19066
rect 9092 19012 9098 19014
rect 9154 19012 9178 19014
rect 9234 19012 9258 19014
rect 9314 19012 9338 19014
rect 9394 19012 9400 19014
rect 9092 19003 9400 19012
rect 10980 18970 11008 21490
rect 14520 21244 14828 21253
rect 14520 21242 14526 21244
rect 14582 21242 14606 21244
rect 14662 21242 14686 21244
rect 14742 21242 14766 21244
rect 14822 21242 14828 21244
rect 14582 21190 14584 21242
rect 14764 21190 14766 21242
rect 14520 21188 14526 21190
rect 14582 21188 14606 21190
rect 14662 21188 14686 21190
rect 14742 21188 14766 21190
rect 14822 21188 14828 21190
rect 14520 21179 14828 21188
rect 15180 20700 15488 20709
rect 15180 20698 15186 20700
rect 15242 20698 15266 20700
rect 15322 20698 15346 20700
rect 15402 20698 15426 20700
rect 15482 20698 15488 20700
rect 15242 20646 15244 20698
rect 15424 20646 15426 20698
rect 15180 20644 15186 20646
rect 15242 20644 15266 20646
rect 15322 20644 15346 20646
rect 15402 20644 15426 20646
rect 15482 20644 15488 20646
rect 15180 20635 15488 20644
rect 14520 20156 14828 20165
rect 14520 20154 14526 20156
rect 14582 20154 14606 20156
rect 14662 20154 14686 20156
rect 14742 20154 14766 20156
rect 14822 20154 14828 20156
rect 14582 20102 14584 20154
rect 14764 20102 14766 20154
rect 14520 20100 14526 20102
rect 14582 20100 14606 20102
rect 14662 20100 14686 20102
rect 14742 20100 14766 20102
rect 14822 20100 14828 20102
rect 14520 20091 14828 20100
rect 15180 19612 15488 19621
rect 15180 19610 15186 19612
rect 15242 19610 15266 19612
rect 15322 19610 15346 19612
rect 15402 19610 15426 19612
rect 15482 19610 15488 19612
rect 15242 19558 15244 19610
rect 15424 19558 15426 19610
rect 15180 19556 15186 19558
rect 15242 19556 15266 19558
rect 15322 19556 15346 19558
rect 15402 19556 15426 19558
rect 15482 19556 15488 19558
rect 15180 19547 15488 19556
rect 14520 19068 14828 19077
rect 14520 19066 14526 19068
rect 14582 19066 14606 19068
rect 14662 19066 14686 19068
rect 14742 19066 14766 19068
rect 14822 19066 14828 19068
rect 14582 19014 14584 19066
rect 14764 19014 14766 19066
rect 14520 19012 14526 19014
rect 14582 19012 14606 19014
rect 14662 19012 14686 19014
rect 14742 19012 14766 19014
rect 14822 19012 14828 19014
rect 14520 19003 14828 19012
rect 4252 18964 4304 18970
rect 4252 18906 4304 18912
rect 10968 18964 11020 18970
rect 10968 18906 11020 18912
rect 4252 18760 4304 18766
rect 4252 18702 4304 18708
rect 10784 18760 10836 18766
rect 10784 18702 10836 18708
rect 4264 18426 4292 18702
rect 4324 18524 4632 18533
rect 4324 18522 4330 18524
rect 4386 18522 4410 18524
rect 4466 18522 4490 18524
rect 4546 18522 4570 18524
rect 4626 18522 4632 18524
rect 4386 18470 4388 18522
rect 4568 18470 4570 18522
rect 4324 18468 4330 18470
rect 4386 18468 4410 18470
rect 4466 18468 4490 18470
rect 4546 18468 4570 18470
rect 4626 18468 4632 18470
rect 4324 18459 4632 18468
rect 9752 18524 10060 18533
rect 9752 18522 9758 18524
rect 9814 18522 9838 18524
rect 9894 18522 9918 18524
rect 9974 18522 9998 18524
rect 10054 18522 10060 18524
rect 9814 18470 9816 18522
rect 9996 18470 9998 18522
rect 9752 18468 9758 18470
rect 9814 18468 9838 18470
rect 9894 18468 9918 18470
rect 9974 18468 9998 18470
rect 10054 18468 10060 18470
rect 9752 18459 10060 18468
rect 10796 18426 10824 18702
rect 15180 18524 15488 18533
rect 15180 18522 15186 18524
rect 15242 18522 15266 18524
rect 15322 18522 15346 18524
rect 15402 18522 15426 18524
rect 15482 18522 15488 18524
rect 15242 18470 15244 18522
rect 15424 18470 15426 18522
rect 15180 18468 15186 18470
rect 15242 18468 15266 18470
rect 15322 18468 15346 18470
rect 15402 18468 15426 18470
rect 15482 18468 15488 18470
rect 15180 18459 15488 18468
rect 4252 18420 4304 18426
rect 4252 18362 4304 18368
rect 10784 18420 10836 18426
rect 10784 18362 10836 18368
rect 4160 18352 4212 18358
rect 4160 18294 4212 18300
rect 1492 18284 1544 18290
rect 1492 18226 1544 18232
rect 1504 17921 1532 18226
rect 4068 18080 4120 18086
rect 4068 18022 4120 18028
rect 3664 17980 3972 17989
rect 3664 17978 3670 17980
rect 3726 17978 3750 17980
rect 3806 17978 3830 17980
rect 3886 17978 3910 17980
rect 3966 17978 3972 17980
rect 3726 17926 3728 17978
rect 3908 17926 3910 17978
rect 3664 17924 3670 17926
rect 3726 17924 3750 17926
rect 3806 17924 3830 17926
rect 3886 17924 3910 17926
rect 3966 17924 3972 17926
rect 1490 17912 1546 17921
rect 3664 17915 3972 17924
rect 1490 17847 1546 17856
rect 3664 16892 3972 16901
rect 3664 16890 3670 16892
rect 3726 16890 3750 16892
rect 3806 16890 3830 16892
rect 3886 16890 3910 16892
rect 3966 16890 3972 16892
rect 3726 16838 3728 16890
rect 3908 16838 3910 16890
rect 3664 16836 3670 16838
rect 3726 16836 3750 16838
rect 3806 16836 3830 16838
rect 3886 16836 3910 16838
rect 3966 16836 3972 16838
rect 3664 16827 3972 16836
rect 3664 15804 3972 15813
rect 3664 15802 3670 15804
rect 3726 15802 3750 15804
rect 3806 15802 3830 15804
rect 3886 15802 3910 15804
rect 3966 15802 3972 15804
rect 3726 15750 3728 15802
rect 3908 15750 3910 15802
rect 3664 15748 3670 15750
rect 3726 15748 3750 15750
rect 3806 15748 3830 15750
rect 3886 15748 3910 15750
rect 3966 15748 3972 15750
rect 3664 15739 3972 15748
rect 3664 14716 3972 14725
rect 3664 14714 3670 14716
rect 3726 14714 3750 14716
rect 3806 14714 3830 14716
rect 3886 14714 3910 14716
rect 3966 14714 3972 14716
rect 3726 14662 3728 14714
rect 3908 14662 3910 14714
rect 3664 14660 3670 14662
rect 3726 14660 3750 14662
rect 3806 14660 3830 14662
rect 3886 14660 3910 14662
rect 3966 14660 3972 14662
rect 3664 14651 3972 14660
rect 3664 13628 3972 13637
rect 3664 13626 3670 13628
rect 3726 13626 3750 13628
rect 3806 13626 3830 13628
rect 3886 13626 3910 13628
rect 3966 13626 3972 13628
rect 3726 13574 3728 13626
rect 3908 13574 3910 13626
rect 3664 13572 3670 13574
rect 3726 13572 3750 13574
rect 3806 13572 3830 13574
rect 3886 13572 3910 13574
rect 3966 13572 3972 13574
rect 3664 13563 3972 13572
rect 3664 12540 3972 12549
rect 3664 12538 3670 12540
rect 3726 12538 3750 12540
rect 3806 12538 3830 12540
rect 3886 12538 3910 12540
rect 3966 12538 3972 12540
rect 3726 12486 3728 12538
rect 3908 12486 3910 12538
rect 3664 12484 3670 12486
rect 3726 12484 3750 12486
rect 3806 12484 3830 12486
rect 3886 12484 3910 12486
rect 3966 12484 3972 12486
rect 3664 12475 3972 12484
rect 3664 11452 3972 11461
rect 3664 11450 3670 11452
rect 3726 11450 3750 11452
rect 3806 11450 3830 11452
rect 3886 11450 3910 11452
rect 3966 11450 3972 11452
rect 3726 11398 3728 11450
rect 3908 11398 3910 11450
rect 3664 11396 3670 11398
rect 3726 11396 3750 11398
rect 3806 11396 3830 11398
rect 3886 11396 3910 11398
rect 3966 11396 3972 11398
rect 3664 11387 3972 11396
rect 3664 10364 3972 10373
rect 3664 10362 3670 10364
rect 3726 10362 3750 10364
rect 3806 10362 3830 10364
rect 3886 10362 3910 10364
rect 3966 10362 3972 10364
rect 3726 10310 3728 10362
rect 3908 10310 3910 10362
rect 3664 10308 3670 10310
rect 3726 10308 3750 10310
rect 3806 10308 3830 10310
rect 3886 10308 3910 10310
rect 3966 10308 3972 10310
rect 3664 10299 3972 10308
rect 3664 9276 3972 9285
rect 3664 9274 3670 9276
rect 3726 9274 3750 9276
rect 3806 9274 3830 9276
rect 3886 9274 3910 9276
rect 3966 9274 3972 9276
rect 3726 9222 3728 9274
rect 3908 9222 3910 9274
rect 3664 9220 3670 9222
rect 3726 9220 3750 9222
rect 3806 9220 3830 9222
rect 3886 9220 3910 9222
rect 3966 9220 3972 9222
rect 3664 9211 3972 9220
rect 4080 8974 4108 18022
rect 4172 9042 4200 18294
rect 15200 18148 15252 18154
rect 15200 18090 15252 18096
rect 9092 17980 9400 17989
rect 9092 17978 9098 17980
rect 9154 17978 9178 17980
rect 9234 17978 9258 17980
rect 9314 17978 9338 17980
rect 9394 17978 9400 17980
rect 9154 17926 9156 17978
rect 9336 17926 9338 17978
rect 9092 17924 9098 17926
rect 9154 17924 9178 17926
rect 9234 17924 9258 17926
rect 9314 17924 9338 17926
rect 9394 17924 9400 17926
rect 9092 17915 9400 17924
rect 14520 17980 14828 17989
rect 14520 17978 14526 17980
rect 14582 17978 14606 17980
rect 14662 17978 14686 17980
rect 14742 17978 14766 17980
rect 14822 17978 14828 17980
rect 14582 17926 14584 17978
rect 14764 17926 14766 17978
rect 14520 17924 14526 17926
rect 14582 17924 14606 17926
rect 14662 17924 14686 17926
rect 14742 17924 14766 17926
rect 14822 17924 14828 17926
rect 14520 17915 14828 17924
rect 15212 17746 15240 18090
rect 17500 18080 17552 18086
rect 17500 18022 17552 18028
rect 17512 17814 17540 18022
rect 18064 17882 18092 21490
rect 19948 21244 20256 21253
rect 19948 21242 19954 21244
rect 20010 21242 20034 21244
rect 20090 21242 20114 21244
rect 20170 21242 20194 21244
rect 20250 21242 20256 21244
rect 20010 21190 20012 21242
rect 20192 21190 20194 21242
rect 19948 21188 19954 21190
rect 20010 21188 20034 21190
rect 20090 21188 20114 21190
rect 20170 21188 20194 21190
rect 20250 21188 20256 21190
rect 19948 21179 20256 21188
rect 20608 20700 20916 20709
rect 20608 20698 20614 20700
rect 20670 20698 20694 20700
rect 20750 20698 20774 20700
rect 20830 20698 20854 20700
rect 20910 20698 20916 20700
rect 20670 20646 20672 20698
rect 20852 20646 20854 20698
rect 20608 20644 20614 20646
rect 20670 20644 20694 20646
rect 20750 20644 20774 20646
rect 20830 20644 20854 20646
rect 20910 20644 20916 20646
rect 20608 20635 20916 20644
rect 19948 20156 20256 20165
rect 19948 20154 19954 20156
rect 20010 20154 20034 20156
rect 20090 20154 20114 20156
rect 20170 20154 20194 20156
rect 20250 20154 20256 20156
rect 20010 20102 20012 20154
rect 20192 20102 20194 20154
rect 19948 20100 19954 20102
rect 20010 20100 20034 20102
rect 20090 20100 20114 20102
rect 20170 20100 20194 20102
rect 20250 20100 20256 20102
rect 19948 20091 20256 20100
rect 22836 19984 22888 19990
rect 22836 19926 22888 19932
rect 22192 19848 22244 19854
rect 22848 19825 22876 19926
rect 22192 19790 22244 19796
rect 22834 19816 22890 19825
rect 20608 19612 20916 19621
rect 20608 19610 20614 19612
rect 20670 19610 20694 19612
rect 20750 19610 20774 19612
rect 20830 19610 20854 19612
rect 20910 19610 20916 19612
rect 20670 19558 20672 19610
rect 20852 19558 20854 19610
rect 20608 19556 20614 19558
rect 20670 19556 20694 19558
rect 20750 19556 20774 19558
rect 20830 19556 20854 19558
rect 20910 19556 20916 19558
rect 20608 19547 20916 19556
rect 19948 19068 20256 19077
rect 19948 19066 19954 19068
rect 20010 19066 20034 19068
rect 20090 19066 20114 19068
rect 20170 19066 20194 19068
rect 20250 19066 20256 19068
rect 20010 19014 20012 19066
rect 20192 19014 20194 19066
rect 19948 19012 19954 19014
rect 20010 19012 20034 19014
rect 20090 19012 20114 19014
rect 20170 19012 20194 19014
rect 20250 19012 20256 19014
rect 19948 19003 20256 19012
rect 20608 18524 20916 18533
rect 20608 18522 20614 18524
rect 20670 18522 20694 18524
rect 20750 18522 20774 18524
rect 20830 18522 20854 18524
rect 20910 18522 20916 18524
rect 20670 18470 20672 18522
rect 20852 18470 20854 18522
rect 20608 18468 20614 18470
rect 20670 18468 20694 18470
rect 20750 18468 20774 18470
rect 20830 18468 20854 18470
rect 20910 18468 20916 18470
rect 20608 18459 20916 18468
rect 22204 18426 22232 19790
rect 22834 19751 22890 19760
rect 22192 18420 22244 18426
rect 22192 18362 22244 18368
rect 18972 18284 19024 18290
rect 18972 18226 19024 18232
rect 18984 17882 19012 18226
rect 19948 17980 20256 17989
rect 19948 17978 19954 17980
rect 20010 17978 20034 17980
rect 20090 17978 20114 17980
rect 20170 17978 20194 17980
rect 20250 17978 20256 17980
rect 20010 17926 20012 17978
rect 20192 17926 20194 17978
rect 19948 17924 19954 17926
rect 20010 17924 20034 17926
rect 20090 17924 20114 17926
rect 20170 17924 20194 17926
rect 20250 17924 20256 17926
rect 19948 17915 20256 17924
rect 18052 17876 18104 17882
rect 18052 17818 18104 17824
rect 18144 17876 18196 17882
rect 18144 17818 18196 17824
rect 18972 17876 19024 17882
rect 18972 17818 19024 17824
rect 17500 17808 17552 17814
rect 17500 17750 17552 17756
rect 15200 17740 15252 17746
rect 15200 17682 15252 17688
rect 17776 17672 17828 17678
rect 17776 17614 17828 17620
rect 4324 17436 4632 17445
rect 4324 17434 4330 17436
rect 4386 17434 4410 17436
rect 4466 17434 4490 17436
rect 4546 17434 4570 17436
rect 4626 17434 4632 17436
rect 4386 17382 4388 17434
rect 4568 17382 4570 17434
rect 4324 17380 4330 17382
rect 4386 17380 4410 17382
rect 4466 17380 4490 17382
rect 4546 17380 4570 17382
rect 4626 17380 4632 17382
rect 4324 17371 4632 17380
rect 9752 17436 10060 17445
rect 9752 17434 9758 17436
rect 9814 17434 9838 17436
rect 9894 17434 9918 17436
rect 9974 17434 9998 17436
rect 10054 17434 10060 17436
rect 9814 17382 9816 17434
rect 9996 17382 9998 17434
rect 9752 17380 9758 17382
rect 9814 17380 9838 17382
rect 9894 17380 9918 17382
rect 9974 17380 9998 17382
rect 10054 17380 10060 17382
rect 9752 17371 10060 17380
rect 15180 17436 15488 17445
rect 15180 17434 15186 17436
rect 15242 17434 15266 17436
rect 15322 17434 15346 17436
rect 15402 17434 15426 17436
rect 15482 17434 15488 17436
rect 15242 17382 15244 17434
rect 15424 17382 15426 17434
rect 15180 17380 15186 17382
rect 15242 17380 15266 17382
rect 15322 17380 15346 17382
rect 15402 17380 15426 17382
rect 15482 17380 15488 17382
rect 15180 17371 15488 17380
rect 9092 16892 9400 16901
rect 9092 16890 9098 16892
rect 9154 16890 9178 16892
rect 9234 16890 9258 16892
rect 9314 16890 9338 16892
rect 9394 16890 9400 16892
rect 9154 16838 9156 16890
rect 9336 16838 9338 16890
rect 9092 16836 9098 16838
rect 9154 16836 9178 16838
rect 9234 16836 9258 16838
rect 9314 16836 9338 16838
rect 9394 16836 9400 16838
rect 9092 16827 9400 16836
rect 14520 16892 14828 16901
rect 14520 16890 14526 16892
rect 14582 16890 14606 16892
rect 14662 16890 14686 16892
rect 14742 16890 14766 16892
rect 14822 16890 14828 16892
rect 14582 16838 14584 16890
rect 14764 16838 14766 16890
rect 14520 16836 14526 16838
rect 14582 16836 14606 16838
rect 14662 16836 14686 16838
rect 14742 16836 14766 16838
rect 14822 16836 14828 16838
rect 14520 16827 14828 16836
rect 4324 16348 4632 16357
rect 4324 16346 4330 16348
rect 4386 16346 4410 16348
rect 4466 16346 4490 16348
rect 4546 16346 4570 16348
rect 4626 16346 4632 16348
rect 4386 16294 4388 16346
rect 4568 16294 4570 16346
rect 4324 16292 4330 16294
rect 4386 16292 4410 16294
rect 4466 16292 4490 16294
rect 4546 16292 4570 16294
rect 4626 16292 4632 16294
rect 4324 16283 4632 16292
rect 9752 16348 10060 16357
rect 9752 16346 9758 16348
rect 9814 16346 9838 16348
rect 9894 16346 9918 16348
rect 9974 16346 9998 16348
rect 10054 16346 10060 16348
rect 9814 16294 9816 16346
rect 9996 16294 9998 16346
rect 9752 16292 9758 16294
rect 9814 16292 9838 16294
rect 9894 16292 9918 16294
rect 9974 16292 9998 16294
rect 10054 16292 10060 16294
rect 9752 16283 10060 16292
rect 15180 16348 15488 16357
rect 15180 16346 15186 16348
rect 15242 16346 15266 16348
rect 15322 16346 15346 16348
rect 15402 16346 15426 16348
rect 15482 16346 15488 16348
rect 15242 16294 15244 16346
rect 15424 16294 15426 16346
rect 15180 16292 15186 16294
rect 15242 16292 15266 16294
rect 15322 16292 15346 16294
rect 15402 16292 15426 16294
rect 15482 16292 15488 16294
rect 15180 16283 15488 16292
rect 9092 15804 9400 15813
rect 9092 15802 9098 15804
rect 9154 15802 9178 15804
rect 9234 15802 9258 15804
rect 9314 15802 9338 15804
rect 9394 15802 9400 15804
rect 9154 15750 9156 15802
rect 9336 15750 9338 15802
rect 9092 15748 9098 15750
rect 9154 15748 9178 15750
rect 9234 15748 9258 15750
rect 9314 15748 9338 15750
rect 9394 15748 9400 15750
rect 9092 15739 9400 15748
rect 14520 15804 14828 15813
rect 14520 15802 14526 15804
rect 14582 15802 14606 15804
rect 14662 15802 14686 15804
rect 14742 15802 14766 15804
rect 14822 15802 14828 15804
rect 14582 15750 14584 15802
rect 14764 15750 14766 15802
rect 14520 15748 14526 15750
rect 14582 15748 14606 15750
rect 14662 15748 14686 15750
rect 14742 15748 14766 15750
rect 14822 15748 14828 15750
rect 14520 15739 14828 15748
rect 4324 15260 4632 15269
rect 4324 15258 4330 15260
rect 4386 15258 4410 15260
rect 4466 15258 4490 15260
rect 4546 15258 4570 15260
rect 4626 15258 4632 15260
rect 4386 15206 4388 15258
rect 4568 15206 4570 15258
rect 4324 15204 4330 15206
rect 4386 15204 4410 15206
rect 4466 15204 4490 15206
rect 4546 15204 4570 15206
rect 4626 15204 4632 15206
rect 4324 15195 4632 15204
rect 9752 15260 10060 15269
rect 9752 15258 9758 15260
rect 9814 15258 9838 15260
rect 9894 15258 9918 15260
rect 9974 15258 9998 15260
rect 10054 15258 10060 15260
rect 9814 15206 9816 15258
rect 9996 15206 9998 15258
rect 9752 15204 9758 15206
rect 9814 15204 9838 15206
rect 9894 15204 9918 15206
rect 9974 15204 9998 15206
rect 10054 15204 10060 15206
rect 9752 15195 10060 15204
rect 15180 15260 15488 15269
rect 15180 15258 15186 15260
rect 15242 15258 15266 15260
rect 15322 15258 15346 15260
rect 15402 15258 15426 15260
rect 15482 15258 15488 15260
rect 15242 15206 15244 15258
rect 15424 15206 15426 15258
rect 15180 15204 15186 15206
rect 15242 15204 15266 15206
rect 15322 15204 15346 15206
rect 15402 15204 15426 15206
rect 15482 15204 15488 15206
rect 15180 15195 15488 15204
rect 9092 14716 9400 14725
rect 9092 14714 9098 14716
rect 9154 14714 9178 14716
rect 9234 14714 9258 14716
rect 9314 14714 9338 14716
rect 9394 14714 9400 14716
rect 9154 14662 9156 14714
rect 9336 14662 9338 14714
rect 9092 14660 9098 14662
rect 9154 14660 9178 14662
rect 9234 14660 9258 14662
rect 9314 14660 9338 14662
rect 9394 14660 9400 14662
rect 9092 14651 9400 14660
rect 14520 14716 14828 14725
rect 14520 14714 14526 14716
rect 14582 14714 14606 14716
rect 14662 14714 14686 14716
rect 14742 14714 14766 14716
rect 14822 14714 14828 14716
rect 14582 14662 14584 14714
rect 14764 14662 14766 14714
rect 14520 14660 14526 14662
rect 14582 14660 14606 14662
rect 14662 14660 14686 14662
rect 14742 14660 14766 14662
rect 14822 14660 14828 14662
rect 14520 14651 14828 14660
rect 4324 14172 4632 14181
rect 4324 14170 4330 14172
rect 4386 14170 4410 14172
rect 4466 14170 4490 14172
rect 4546 14170 4570 14172
rect 4626 14170 4632 14172
rect 4386 14118 4388 14170
rect 4568 14118 4570 14170
rect 4324 14116 4330 14118
rect 4386 14116 4410 14118
rect 4466 14116 4490 14118
rect 4546 14116 4570 14118
rect 4626 14116 4632 14118
rect 4324 14107 4632 14116
rect 9752 14172 10060 14181
rect 9752 14170 9758 14172
rect 9814 14170 9838 14172
rect 9894 14170 9918 14172
rect 9974 14170 9998 14172
rect 10054 14170 10060 14172
rect 9814 14118 9816 14170
rect 9996 14118 9998 14170
rect 9752 14116 9758 14118
rect 9814 14116 9838 14118
rect 9894 14116 9918 14118
rect 9974 14116 9998 14118
rect 10054 14116 10060 14118
rect 9752 14107 10060 14116
rect 15180 14172 15488 14181
rect 15180 14170 15186 14172
rect 15242 14170 15266 14172
rect 15322 14170 15346 14172
rect 15402 14170 15426 14172
rect 15482 14170 15488 14172
rect 15242 14118 15244 14170
rect 15424 14118 15426 14170
rect 15180 14116 15186 14118
rect 15242 14116 15266 14118
rect 15322 14116 15346 14118
rect 15402 14116 15426 14118
rect 15482 14116 15488 14118
rect 15180 14107 15488 14116
rect 9092 13628 9400 13637
rect 9092 13626 9098 13628
rect 9154 13626 9178 13628
rect 9234 13626 9258 13628
rect 9314 13626 9338 13628
rect 9394 13626 9400 13628
rect 9154 13574 9156 13626
rect 9336 13574 9338 13626
rect 9092 13572 9098 13574
rect 9154 13572 9178 13574
rect 9234 13572 9258 13574
rect 9314 13572 9338 13574
rect 9394 13572 9400 13574
rect 9092 13563 9400 13572
rect 14520 13628 14828 13637
rect 14520 13626 14526 13628
rect 14582 13626 14606 13628
rect 14662 13626 14686 13628
rect 14742 13626 14766 13628
rect 14822 13626 14828 13628
rect 14582 13574 14584 13626
rect 14764 13574 14766 13626
rect 14520 13572 14526 13574
rect 14582 13572 14606 13574
rect 14662 13572 14686 13574
rect 14742 13572 14766 13574
rect 14822 13572 14828 13574
rect 14520 13563 14828 13572
rect 4324 13084 4632 13093
rect 4324 13082 4330 13084
rect 4386 13082 4410 13084
rect 4466 13082 4490 13084
rect 4546 13082 4570 13084
rect 4626 13082 4632 13084
rect 4386 13030 4388 13082
rect 4568 13030 4570 13082
rect 4324 13028 4330 13030
rect 4386 13028 4410 13030
rect 4466 13028 4490 13030
rect 4546 13028 4570 13030
rect 4626 13028 4632 13030
rect 4324 13019 4632 13028
rect 9752 13084 10060 13093
rect 9752 13082 9758 13084
rect 9814 13082 9838 13084
rect 9894 13082 9918 13084
rect 9974 13082 9998 13084
rect 10054 13082 10060 13084
rect 9814 13030 9816 13082
rect 9996 13030 9998 13082
rect 9752 13028 9758 13030
rect 9814 13028 9838 13030
rect 9894 13028 9918 13030
rect 9974 13028 9998 13030
rect 10054 13028 10060 13030
rect 9752 13019 10060 13028
rect 15180 13084 15488 13093
rect 15180 13082 15186 13084
rect 15242 13082 15266 13084
rect 15322 13082 15346 13084
rect 15402 13082 15426 13084
rect 15482 13082 15488 13084
rect 15242 13030 15244 13082
rect 15424 13030 15426 13082
rect 15180 13028 15186 13030
rect 15242 13028 15266 13030
rect 15322 13028 15346 13030
rect 15402 13028 15426 13030
rect 15482 13028 15488 13030
rect 15180 13019 15488 13028
rect 9092 12540 9400 12549
rect 9092 12538 9098 12540
rect 9154 12538 9178 12540
rect 9234 12538 9258 12540
rect 9314 12538 9338 12540
rect 9394 12538 9400 12540
rect 9154 12486 9156 12538
rect 9336 12486 9338 12538
rect 9092 12484 9098 12486
rect 9154 12484 9178 12486
rect 9234 12484 9258 12486
rect 9314 12484 9338 12486
rect 9394 12484 9400 12486
rect 9092 12475 9400 12484
rect 14520 12540 14828 12549
rect 14520 12538 14526 12540
rect 14582 12538 14606 12540
rect 14662 12538 14686 12540
rect 14742 12538 14766 12540
rect 14822 12538 14828 12540
rect 14582 12486 14584 12538
rect 14764 12486 14766 12538
rect 14520 12484 14526 12486
rect 14582 12484 14606 12486
rect 14662 12484 14686 12486
rect 14742 12484 14766 12486
rect 14822 12484 14828 12486
rect 14520 12475 14828 12484
rect 4324 11996 4632 12005
rect 4324 11994 4330 11996
rect 4386 11994 4410 11996
rect 4466 11994 4490 11996
rect 4546 11994 4570 11996
rect 4626 11994 4632 11996
rect 4386 11942 4388 11994
rect 4568 11942 4570 11994
rect 4324 11940 4330 11942
rect 4386 11940 4410 11942
rect 4466 11940 4490 11942
rect 4546 11940 4570 11942
rect 4626 11940 4632 11942
rect 4324 11931 4632 11940
rect 9752 11996 10060 12005
rect 9752 11994 9758 11996
rect 9814 11994 9838 11996
rect 9894 11994 9918 11996
rect 9974 11994 9998 11996
rect 10054 11994 10060 11996
rect 9814 11942 9816 11994
rect 9996 11942 9998 11994
rect 9752 11940 9758 11942
rect 9814 11940 9838 11942
rect 9894 11940 9918 11942
rect 9974 11940 9998 11942
rect 10054 11940 10060 11942
rect 9752 11931 10060 11940
rect 15180 11996 15488 12005
rect 15180 11994 15186 11996
rect 15242 11994 15266 11996
rect 15322 11994 15346 11996
rect 15402 11994 15426 11996
rect 15482 11994 15488 11996
rect 15242 11942 15244 11994
rect 15424 11942 15426 11994
rect 15180 11940 15186 11942
rect 15242 11940 15266 11942
rect 15322 11940 15346 11942
rect 15402 11940 15426 11942
rect 15482 11940 15488 11942
rect 15180 11931 15488 11940
rect 9092 11452 9400 11461
rect 9092 11450 9098 11452
rect 9154 11450 9178 11452
rect 9234 11450 9258 11452
rect 9314 11450 9338 11452
rect 9394 11450 9400 11452
rect 9154 11398 9156 11450
rect 9336 11398 9338 11450
rect 9092 11396 9098 11398
rect 9154 11396 9178 11398
rect 9234 11396 9258 11398
rect 9314 11396 9338 11398
rect 9394 11396 9400 11398
rect 9092 11387 9400 11396
rect 14520 11452 14828 11461
rect 14520 11450 14526 11452
rect 14582 11450 14606 11452
rect 14662 11450 14686 11452
rect 14742 11450 14766 11452
rect 14822 11450 14828 11452
rect 14582 11398 14584 11450
rect 14764 11398 14766 11450
rect 14520 11396 14526 11398
rect 14582 11396 14606 11398
rect 14662 11396 14686 11398
rect 14742 11396 14766 11398
rect 14822 11396 14828 11398
rect 14520 11387 14828 11396
rect 4324 10908 4632 10917
rect 4324 10906 4330 10908
rect 4386 10906 4410 10908
rect 4466 10906 4490 10908
rect 4546 10906 4570 10908
rect 4626 10906 4632 10908
rect 4386 10854 4388 10906
rect 4568 10854 4570 10906
rect 4324 10852 4330 10854
rect 4386 10852 4410 10854
rect 4466 10852 4490 10854
rect 4546 10852 4570 10854
rect 4626 10852 4632 10854
rect 4324 10843 4632 10852
rect 9752 10908 10060 10917
rect 9752 10906 9758 10908
rect 9814 10906 9838 10908
rect 9894 10906 9918 10908
rect 9974 10906 9998 10908
rect 10054 10906 10060 10908
rect 9814 10854 9816 10906
rect 9996 10854 9998 10906
rect 9752 10852 9758 10854
rect 9814 10852 9838 10854
rect 9894 10852 9918 10854
rect 9974 10852 9998 10854
rect 10054 10852 10060 10854
rect 9752 10843 10060 10852
rect 15180 10908 15488 10917
rect 15180 10906 15186 10908
rect 15242 10906 15266 10908
rect 15322 10906 15346 10908
rect 15402 10906 15426 10908
rect 15482 10906 15488 10908
rect 15242 10854 15244 10906
rect 15424 10854 15426 10906
rect 15180 10852 15186 10854
rect 15242 10852 15266 10854
rect 15322 10852 15346 10854
rect 15402 10852 15426 10854
rect 15482 10852 15488 10854
rect 15180 10843 15488 10852
rect 9092 10364 9400 10373
rect 9092 10362 9098 10364
rect 9154 10362 9178 10364
rect 9234 10362 9258 10364
rect 9314 10362 9338 10364
rect 9394 10362 9400 10364
rect 9154 10310 9156 10362
rect 9336 10310 9338 10362
rect 9092 10308 9098 10310
rect 9154 10308 9178 10310
rect 9234 10308 9258 10310
rect 9314 10308 9338 10310
rect 9394 10308 9400 10310
rect 9092 10299 9400 10308
rect 14520 10364 14828 10373
rect 14520 10362 14526 10364
rect 14582 10362 14606 10364
rect 14662 10362 14686 10364
rect 14742 10362 14766 10364
rect 14822 10362 14828 10364
rect 14582 10310 14584 10362
rect 14764 10310 14766 10362
rect 14520 10308 14526 10310
rect 14582 10308 14606 10310
rect 14662 10308 14686 10310
rect 14742 10308 14766 10310
rect 14822 10308 14828 10310
rect 14520 10299 14828 10308
rect 17788 9994 17816 17614
rect 18156 10266 18184 17818
rect 18236 17536 18288 17542
rect 18236 17478 18288 17484
rect 18144 10260 18196 10266
rect 18144 10202 18196 10208
rect 16856 9988 16908 9994
rect 16856 9930 16908 9936
rect 17776 9988 17828 9994
rect 17776 9930 17828 9936
rect 4324 9820 4632 9829
rect 4324 9818 4330 9820
rect 4386 9818 4410 9820
rect 4466 9818 4490 9820
rect 4546 9818 4570 9820
rect 4626 9818 4632 9820
rect 4386 9766 4388 9818
rect 4568 9766 4570 9818
rect 4324 9764 4330 9766
rect 4386 9764 4410 9766
rect 4466 9764 4490 9766
rect 4546 9764 4570 9766
rect 4626 9764 4632 9766
rect 4324 9755 4632 9764
rect 9752 9820 10060 9829
rect 9752 9818 9758 9820
rect 9814 9818 9838 9820
rect 9894 9818 9918 9820
rect 9974 9818 9998 9820
rect 10054 9818 10060 9820
rect 9814 9766 9816 9818
rect 9996 9766 9998 9818
rect 9752 9764 9758 9766
rect 9814 9764 9838 9766
rect 9894 9764 9918 9766
rect 9974 9764 9998 9766
rect 10054 9764 10060 9766
rect 9752 9755 10060 9764
rect 15180 9820 15488 9829
rect 15180 9818 15186 9820
rect 15242 9818 15266 9820
rect 15322 9818 15346 9820
rect 15402 9818 15426 9820
rect 15482 9818 15488 9820
rect 15242 9766 15244 9818
rect 15424 9766 15426 9818
rect 15180 9764 15186 9766
rect 15242 9764 15266 9766
rect 15322 9764 15346 9766
rect 15402 9764 15426 9766
rect 15482 9764 15488 9766
rect 15180 9755 15488 9764
rect 9092 9276 9400 9285
rect 9092 9274 9098 9276
rect 9154 9274 9178 9276
rect 9234 9274 9258 9276
rect 9314 9274 9338 9276
rect 9394 9274 9400 9276
rect 9154 9222 9156 9274
rect 9336 9222 9338 9274
rect 9092 9220 9098 9222
rect 9154 9220 9178 9222
rect 9234 9220 9258 9222
rect 9314 9220 9338 9222
rect 9394 9220 9400 9222
rect 9092 9211 9400 9220
rect 14520 9276 14828 9285
rect 14520 9274 14526 9276
rect 14582 9274 14606 9276
rect 14662 9274 14686 9276
rect 14742 9274 14766 9276
rect 14822 9274 14828 9276
rect 14582 9222 14584 9274
rect 14764 9222 14766 9274
rect 14520 9220 14526 9222
rect 14582 9220 14606 9222
rect 14662 9220 14686 9222
rect 14742 9220 14766 9222
rect 14822 9220 14828 9222
rect 14520 9211 14828 9220
rect 4160 9036 4212 9042
rect 4160 8978 4212 8984
rect 4712 9036 4764 9042
rect 4712 8978 4764 8984
rect 4068 8968 4120 8974
rect 938 8936 994 8945
rect 4068 8910 4120 8916
rect 938 8871 940 8880
rect 992 8871 994 8880
rect 940 8842 992 8848
rect 3664 8188 3972 8197
rect 3664 8186 3670 8188
rect 3726 8186 3750 8188
rect 3806 8186 3830 8188
rect 3886 8186 3910 8188
rect 3966 8186 3972 8188
rect 3726 8134 3728 8186
rect 3908 8134 3910 8186
rect 3664 8132 3670 8134
rect 3726 8132 3750 8134
rect 3806 8132 3830 8134
rect 3886 8132 3910 8134
rect 3966 8132 3972 8134
rect 3664 8123 3972 8132
rect 3664 7100 3972 7109
rect 3664 7098 3670 7100
rect 3726 7098 3750 7100
rect 3806 7098 3830 7100
rect 3886 7098 3910 7100
rect 3966 7098 3972 7100
rect 3726 7046 3728 7098
rect 3908 7046 3910 7098
rect 3664 7044 3670 7046
rect 3726 7044 3750 7046
rect 3806 7044 3830 7046
rect 3886 7044 3910 7046
rect 3966 7044 3972 7046
rect 3664 7035 3972 7044
rect 3664 6012 3972 6021
rect 3664 6010 3670 6012
rect 3726 6010 3750 6012
rect 3806 6010 3830 6012
rect 3886 6010 3910 6012
rect 3966 6010 3972 6012
rect 3726 5958 3728 6010
rect 3908 5958 3910 6010
rect 3664 5956 3670 5958
rect 3726 5956 3750 5958
rect 3806 5956 3830 5958
rect 3886 5956 3910 5958
rect 3966 5956 3972 5958
rect 3664 5947 3972 5956
rect 3664 4924 3972 4933
rect 3664 4922 3670 4924
rect 3726 4922 3750 4924
rect 3806 4922 3830 4924
rect 3886 4922 3910 4924
rect 3966 4922 3972 4924
rect 3726 4870 3728 4922
rect 3908 4870 3910 4922
rect 3664 4868 3670 4870
rect 3726 4868 3750 4870
rect 3806 4868 3830 4870
rect 3886 4868 3910 4870
rect 3966 4868 3972 4870
rect 3664 4859 3972 4868
rect 4080 4146 4108 8910
rect 4324 8732 4632 8741
rect 4324 8730 4330 8732
rect 4386 8730 4410 8732
rect 4466 8730 4490 8732
rect 4546 8730 4570 8732
rect 4626 8730 4632 8732
rect 4386 8678 4388 8730
rect 4568 8678 4570 8730
rect 4324 8676 4330 8678
rect 4386 8676 4410 8678
rect 4466 8676 4490 8678
rect 4546 8676 4570 8678
rect 4626 8676 4632 8678
rect 4324 8667 4632 8676
rect 4324 7644 4632 7653
rect 4324 7642 4330 7644
rect 4386 7642 4410 7644
rect 4466 7642 4490 7644
rect 4546 7642 4570 7644
rect 4626 7642 4632 7644
rect 4386 7590 4388 7642
rect 4568 7590 4570 7642
rect 4324 7588 4330 7590
rect 4386 7588 4410 7590
rect 4466 7588 4490 7590
rect 4546 7588 4570 7590
rect 4626 7588 4632 7590
rect 4324 7579 4632 7588
rect 4324 6556 4632 6565
rect 4324 6554 4330 6556
rect 4386 6554 4410 6556
rect 4466 6554 4490 6556
rect 4546 6554 4570 6556
rect 4626 6554 4632 6556
rect 4386 6502 4388 6554
rect 4568 6502 4570 6554
rect 4324 6500 4330 6502
rect 4386 6500 4410 6502
rect 4466 6500 4490 6502
rect 4546 6500 4570 6502
rect 4626 6500 4632 6502
rect 4324 6491 4632 6500
rect 4324 5468 4632 5477
rect 4324 5466 4330 5468
rect 4386 5466 4410 5468
rect 4466 5466 4490 5468
rect 4546 5466 4570 5468
rect 4626 5466 4632 5468
rect 4386 5414 4388 5466
rect 4568 5414 4570 5466
rect 4324 5412 4330 5414
rect 4386 5412 4410 5414
rect 4466 5412 4490 5414
rect 4546 5412 4570 5414
rect 4626 5412 4632 5414
rect 4324 5403 4632 5412
rect 4324 4380 4632 4389
rect 4324 4378 4330 4380
rect 4386 4378 4410 4380
rect 4466 4378 4490 4380
rect 4546 4378 4570 4380
rect 4626 4378 4632 4380
rect 4386 4326 4388 4378
rect 4568 4326 4570 4378
rect 4324 4324 4330 4326
rect 4386 4324 4410 4326
rect 4466 4324 4490 4326
rect 4546 4324 4570 4326
rect 4626 4324 4632 4326
rect 4324 4315 4632 4324
rect 4724 4146 4752 8978
rect 8024 8968 8076 8974
rect 8024 8910 8076 8916
rect 8036 4146 8064 8910
rect 9752 8732 10060 8741
rect 9752 8730 9758 8732
rect 9814 8730 9838 8732
rect 9894 8730 9918 8732
rect 9974 8730 9998 8732
rect 10054 8730 10060 8732
rect 9814 8678 9816 8730
rect 9996 8678 9998 8730
rect 9752 8676 9758 8678
rect 9814 8676 9838 8678
rect 9894 8676 9918 8678
rect 9974 8676 9998 8678
rect 10054 8676 10060 8678
rect 9752 8667 10060 8676
rect 15180 8732 15488 8741
rect 15180 8730 15186 8732
rect 15242 8730 15266 8732
rect 15322 8730 15346 8732
rect 15402 8730 15426 8732
rect 15482 8730 15488 8732
rect 15242 8678 15244 8730
rect 15424 8678 15426 8730
rect 15180 8676 15186 8678
rect 15242 8676 15266 8678
rect 15322 8676 15346 8678
rect 15402 8676 15426 8678
rect 15482 8676 15488 8678
rect 15180 8667 15488 8676
rect 9092 8188 9400 8197
rect 9092 8186 9098 8188
rect 9154 8186 9178 8188
rect 9234 8186 9258 8188
rect 9314 8186 9338 8188
rect 9394 8186 9400 8188
rect 9154 8134 9156 8186
rect 9336 8134 9338 8186
rect 9092 8132 9098 8134
rect 9154 8132 9178 8134
rect 9234 8132 9258 8134
rect 9314 8132 9338 8134
rect 9394 8132 9400 8134
rect 9092 8123 9400 8132
rect 14520 8188 14828 8197
rect 14520 8186 14526 8188
rect 14582 8186 14606 8188
rect 14662 8186 14686 8188
rect 14742 8186 14766 8188
rect 14822 8186 14828 8188
rect 14582 8134 14584 8186
rect 14764 8134 14766 8186
rect 14520 8132 14526 8134
rect 14582 8132 14606 8134
rect 14662 8132 14686 8134
rect 14742 8132 14766 8134
rect 14822 8132 14828 8134
rect 14520 8123 14828 8132
rect 9752 7644 10060 7653
rect 9752 7642 9758 7644
rect 9814 7642 9838 7644
rect 9894 7642 9918 7644
rect 9974 7642 9998 7644
rect 10054 7642 10060 7644
rect 9814 7590 9816 7642
rect 9996 7590 9998 7642
rect 9752 7588 9758 7590
rect 9814 7588 9838 7590
rect 9894 7588 9918 7590
rect 9974 7588 9998 7590
rect 10054 7588 10060 7590
rect 9752 7579 10060 7588
rect 15180 7644 15488 7653
rect 15180 7642 15186 7644
rect 15242 7642 15266 7644
rect 15322 7642 15346 7644
rect 15402 7642 15426 7644
rect 15482 7642 15488 7644
rect 15242 7590 15244 7642
rect 15424 7590 15426 7642
rect 15180 7588 15186 7590
rect 15242 7588 15266 7590
rect 15322 7588 15346 7590
rect 15402 7588 15426 7590
rect 15482 7588 15488 7590
rect 15180 7579 15488 7588
rect 9092 7100 9400 7109
rect 9092 7098 9098 7100
rect 9154 7098 9178 7100
rect 9234 7098 9258 7100
rect 9314 7098 9338 7100
rect 9394 7098 9400 7100
rect 9154 7046 9156 7098
rect 9336 7046 9338 7098
rect 9092 7044 9098 7046
rect 9154 7044 9178 7046
rect 9234 7044 9258 7046
rect 9314 7044 9338 7046
rect 9394 7044 9400 7046
rect 9092 7035 9400 7044
rect 14520 7100 14828 7109
rect 14520 7098 14526 7100
rect 14582 7098 14606 7100
rect 14662 7098 14686 7100
rect 14742 7098 14766 7100
rect 14822 7098 14828 7100
rect 14582 7046 14584 7098
rect 14764 7046 14766 7098
rect 14520 7044 14526 7046
rect 14582 7044 14606 7046
rect 14662 7044 14686 7046
rect 14742 7044 14766 7046
rect 14822 7044 14828 7046
rect 14520 7035 14828 7044
rect 9752 6556 10060 6565
rect 9752 6554 9758 6556
rect 9814 6554 9838 6556
rect 9894 6554 9918 6556
rect 9974 6554 9998 6556
rect 10054 6554 10060 6556
rect 9814 6502 9816 6554
rect 9996 6502 9998 6554
rect 9752 6500 9758 6502
rect 9814 6500 9838 6502
rect 9894 6500 9918 6502
rect 9974 6500 9998 6502
rect 10054 6500 10060 6502
rect 9752 6491 10060 6500
rect 15180 6556 15488 6565
rect 15180 6554 15186 6556
rect 15242 6554 15266 6556
rect 15322 6554 15346 6556
rect 15402 6554 15426 6556
rect 15482 6554 15488 6556
rect 15242 6502 15244 6554
rect 15424 6502 15426 6554
rect 15180 6500 15186 6502
rect 15242 6500 15266 6502
rect 15322 6500 15346 6502
rect 15402 6500 15426 6502
rect 15482 6500 15488 6502
rect 15180 6491 15488 6500
rect 9092 6012 9400 6021
rect 9092 6010 9098 6012
rect 9154 6010 9178 6012
rect 9234 6010 9258 6012
rect 9314 6010 9338 6012
rect 9394 6010 9400 6012
rect 9154 5958 9156 6010
rect 9336 5958 9338 6010
rect 9092 5956 9098 5958
rect 9154 5956 9178 5958
rect 9234 5956 9258 5958
rect 9314 5956 9338 5958
rect 9394 5956 9400 5958
rect 9092 5947 9400 5956
rect 14520 6012 14828 6021
rect 14520 6010 14526 6012
rect 14582 6010 14606 6012
rect 14662 6010 14686 6012
rect 14742 6010 14766 6012
rect 14822 6010 14828 6012
rect 14582 5958 14584 6010
rect 14764 5958 14766 6010
rect 14520 5956 14526 5958
rect 14582 5956 14606 5958
rect 14662 5956 14686 5958
rect 14742 5956 14766 5958
rect 14822 5956 14828 5958
rect 14520 5947 14828 5956
rect 9752 5468 10060 5477
rect 9752 5466 9758 5468
rect 9814 5466 9838 5468
rect 9894 5466 9918 5468
rect 9974 5466 9998 5468
rect 10054 5466 10060 5468
rect 9814 5414 9816 5466
rect 9996 5414 9998 5466
rect 9752 5412 9758 5414
rect 9814 5412 9838 5414
rect 9894 5412 9918 5414
rect 9974 5412 9998 5414
rect 10054 5412 10060 5414
rect 9752 5403 10060 5412
rect 15180 5468 15488 5477
rect 15180 5466 15186 5468
rect 15242 5466 15266 5468
rect 15322 5466 15346 5468
rect 15402 5466 15426 5468
rect 15482 5466 15488 5468
rect 15242 5414 15244 5466
rect 15424 5414 15426 5466
rect 15180 5412 15186 5414
rect 15242 5412 15266 5414
rect 15322 5412 15346 5414
rect 15402 5412 15426 5414
rect 15482 5412 15488 5414
rect 15180 5403 15488 5412
rect 16868 5234 16896 9930
rect 16856 5228 16908 5234
rect 16856 5170 16908 5176
rect 9092 4924 9400 4933
rect 9092 4922 9098 4924
rect 9154 4922 9178 4924
rect 9234 4922 9258 4924
rect 9314 4922 9338 4924
rect 9394 4922 9400 4924
rect 9154 4870 9156 4922
rect 9336 4870 9338 4922
rect 9092 4868 9098 4870
rect 9154 4868 9178 4870
rect 9234 4868 9258 4870
rect 9314 4868 9338 4870
rect 9394 4868 9400 4870
rect 9092 4859 9400 4868
rect 14520 4924 14828 4933
rect 14520 4922 14526 4924
rect 14582 4922 14606 4924
rect 14662 4922 14686 4924
rect 14742 4922 14766 4924
rect 14822 4922 14828 4924
rect 14582 4870 14584 4922
rect 14764 4870 14766 4922
rect 14520 4868 14526 4870
rect 14582 4868 14606 4870
rect 14662 4868 14686 4870
rect 14742 4868 14766 4870
rect 14822 4868 14828 4870
rect 14520 4859 14828 4868
rect 9752 4380 10060 4389
rect 9752 4378 9758 4380
rect 9814 4378 9838 4380
rect 9894 4378 9918 4380
rect 9974 4378 9998 4380
rect 10054 4378 10060 4380
rect 9814 4326 9816 4378
rect 9996 4326 9998 4378
rect 9752 4324 9758 4326
rect 9814 4324 9838 4326
rect 9894 4324 9918 4326
rect 9974 4324 9998 4326
rect 10054 4324 10060 4326
rect 9752 4315 10060 4324
rect 15180 4380 15488 4389
rect 15180 4378 15186 4380
rect 15242 4378 15266 4380
rect 15322 4378 15346 4380
rect 15402 4378 15426 4380
rect 15482 4378 15488 4380
rect 15242 4326 15244 4378
rect 15424 4326 15426 4378
rect 15180 4324 15186 4326
rect 15242 4324 15266 4326
rect 15322 4324 15346 4326
rect 15402 4324 15426 4326
rect 15482 4324 15488 4326
rect 15180 4315 15488 4324
rect 8220 4146 8432 4162
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 4712 4140 4764 4146
rect 4712 4082 4764 4088
rect 8024 4140 8076 4146
rect 8024 4082 8076 4088
rect 8208 4140 8444 4146
rect 8260 4134 8392 4140
rect 8208 4082 8260 4088
rect 8392 4082 8444 4088
rect 3664 3836 3972 3845
rect 3664 3834 3670 3836
rect 3726 3834 3750 3836
rect 3806 3834 3830 3836
rect 3886 3834 3910 3836
rect 3966 3834 3972 3836
rect 3726 3782 3728 3834
rect 3908 3782 3910 3834
rect 3664 3780 3670 3782
rect 3726 3780 3750 3782
rect 3806 3780 3830 3782
rect 3886 3780 3910 3782
rect 3966 3780 3972 3782
rect 3664 3771 3972 3780
rect 4324 3292 4632 3301
rect 4324 3290 4330 3292
rect 4386 3290 4410 3292
rect 4466 3290 4490 3292
rect 4546 3290 4570 3292
rect 4626 3290 4632 3292
rect 4386 3238 4388 3290
rect 4568 3238 4570 3290
rect 4324 3236 4330 3238
rect 4386 3236 4410 3238
rect 4466 3236 4490 3238
rect 4546 3236 4570 3238
rect 4626 3236 4632 3238
rect 4324 3227 4632 3236
rect 3664 2748 3972 2757
rect 3664 2746 3670 2748
rect 3726 2746 3750 2748
rect 3806 2746 3830 2748
rect 3886 2746 3910 2748
rect 3966 2746 3972 2748
rect 3726 2694 3728 2746
rect 3908 2694 3910 2746
rect 3664 2692 3670 2694
rect 3726 2692 3750 2694
rect 3806 2692 3830 2694
rect 3886 2692 3910 2694
rect 3966 2692 3972 2694
rect 3664 2683 3972 2692
rect 4724 2650 4752 4082
rect 16868 4078 16896 5170
rect 16948 5160 17000 5166
rect 16948 5102 17000 5108
rect 16960 4146 16988 5102
rect 17132 5024 17184 5030
rect 17132 4966 17184 4972
rect 16948 4140 17000 4146
rect 16948 4082 17000 4088
rect 16856 4072 16908 4078
rect 16856 4014 16908 4020
rect 8484 3936 8536 3942
rect 8484 3878 8536 3884
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 8496 2446 8524 3878
rect 9092 3836 9400 3845
rect 9092 3834 9098 3836
rect 9154 3834 9178 3836
rect 9234 3834 9258 3836
rect 9314 3834 9338 3836
rect 9394 3834 9400 3836
rect 9154 3782 9156 3834
rect 9336 3782 9338 3834
rect 9092 3780 9098 3782
rect 9154 3780 9178 3782
rect 9234 3780 9258 3782
rect 9314 3780 9338 3782
rect 9394 3780 9400 3782
rect 9092 3771 9400 3780
rect 14520 3836 14828 3845
rect 14520 3834 14526 3836
rect 14582 3834 14606 3836
rect 14662 3834 14686 3836
rect 14742 3834 14766 3836
rect 14822 3834 14828 3836
rect 14582 3782 14584 3834
rect 14764 3782 14766 3834
rect 14520 3780 14526 3782
rect 14582 3780 14606 3782
rect 14662 3780 14686 3782
rect 14742 3780 14766 3782
rect 14822 3780 14828 3782
rect 14520 3771 14828 3780
rect 9752 3292 10060 3301
rect 9752 3290 9758 3292
rect 9814 3290 9838 3292
rect 9894 3290 9918 3292
rect 9974 3290 9998 3292
rect 10054 3290 10060 3292
rect 9814 3238 9816 3290
rect 9996 3238 9998 3290
rect 9752 3236 9758 3238
rect 9814 3236 9838 3238
rect 9894 3236 9918 3238
rect 9974 3236 9998 3238
rect 10054 3236 10060 3238
rect 9752 3227 10060 3236
rect 15180 3292 15488 3301
rect 15180 3290 15186 3292
rect 15242 3290 15266 3292
rect 15322 3290 15346 3292
rect 15402 3290 15426 3292
rect 15482 3290 15488 3292
rect 15242 3238 15244 3290
rect 15424 3238 15426 3290
rect 15180 3236 15186 3238
rect 15242 3236 15266 3238
rect 15322 3236 15346 3238
rect 15402 3236 15426 3238
rect 15482 3236 15488 3238
rect 15180 3227 15488 3236
rect 9092 2748 9400 2757
rect 9092 2746 9098 2748
rect 9154 2746 9178 2748
rect 9234 2746 9258 2748
rect 9314 2746 9338 2748
rect 9394 2746 9400 2748
rect 9154 2694 9156 2746
rect 9336 2694 9338 2746
rect 9092 2692 9098 2694
rect 9154 2692 9178 2694
rect 9234 2692 9258 2694
rect 9314 2692 9338 2694
rect 9394 2692 9400 2694
rect 9092 2683 9400 2692
rect 14520 2748 14828 2757
rect 14520 2746 14526 2748
rect 14582 2746 14606 2748
rect 14662 2746 14686 2748
rect 14742 2746 14766 2748
rect 14822 2746 14828 2748
rect 14582 2694 14584 2746
rect 14764 2694 14766 2746
rect 14520 2692 14526 2694
rect 14582 2692 14606 2694
rect 14662 2692 14686 2694
rect 14742 2692 14766 2694
rect 14822 2692 14828 2694
rect 14520 2683 14828 2692
rect 17144 2446 17172 4966
rect 18156 4214 18184 10202
rect 18248 10062 18276 17478
rect 20608 17436 20916 17445
rect 20608 17434 20614 17436
rect 20670 17434 20694 17436
rect 20750 17434 20774 17436
rect 20830 17434 20854 17436
rect 20910 17434 20916 17436
rect 20670 17382 20672 17434
rect 20852 17382 20854 17434
rect 20608 17380 20614 17382
rect 20670 17380 20694 17382
rect 20750 17380 20774 17382
rect 20830 17380 20854 17382
rect 20910 17380 20916 17382
rect 20608 17371 20916 17380
rect 19948 16892 20256 16901
rect 19948 16890 19954 16892
rect 20010 16890 20034 16892
rect 20090 16890 20114 16892
rect 20170 16890 20194 16892
rect 20250 16890 20256 16892
rect 20010 16838 20012 16890
rect 20192 16838 20194 16890
rect 19948 16836 19954 16838
rect 20010 16836 20034 16838
rect 20090 16836 20114 16838
rect 20170 16836 20194 16838
rect 20250 16836 20256 16838
rect 19948 16827 20256 16836
rect 20608 16348 20916 16357
rect 20608 16346 20614 16348
rect 20670 16346 20694 16348
rect 20750 16346 20774 16348
rect 20830 16346 20854 16348
rect 20910 16346 20916 16348
rect 20670 16294 20672 16346
rect 20852 16294 20854 16346
rect 20608 16292 20614 16294
rect 20670 16292 20694 16294
rect 20750 16292 20774 16294
rect 20830 16292 20854 16294
rect 20910 16292 20916 16294
rect 20608 16283 20916 16292
rect 19948 15804 20256 15813
rect 19948 15802 19954 15804
rect 20010 15802 20034 15804
rect 20090 15802 20114 15804
rect 20170 15802 20194 15804
rect 20250 15802 20256 15804
rect 20010 15750 20012 15802
rect 20192 15750 20194 15802
rect 19948 15748 19954 15750
rect 20010 15748 20034 15750
rect 20090 15748 20114 15750
rect 20170 15748 20194 15750
rect 20250 15748 20256 15750
rect 19948 15739 20256 15748
rect 20608 15260 20916 15269
rect 20608 15258 20614 15260
rect 20670 15258 20694 15260
rect 20750 15258 20774 15260
rect 20830 15258 20854 15260
rect 20910 15258 20916 15260
rect 20670 15206 20672 15258
rect 20852 15206 20854 15258
rect 20608 15204 20614 15206
rect 20670 15204 20694 15206
rect 20750 15204 20774 15206
rect 20830 15204 20854 15206
rect 20910 15204 20916 15206
rect 20608 15195 20916 15204
rect 19948 14716 20256 14725
rect 19948 14714 19954 14716
rect 20010 14714 20034 14716
rect 20090 14714 20114 14716
rect 20170 14714 20194 14716
rect 20250 14714 20256 14716
rect 20010 14662 20012 14714
rect 20192 14662 20194 14714
rect 19948 14660 19954 14662
rect 20010 14660 20034 14662
rect 20090 14660 20114 14662
rect 20170 14660 20194 14662
rect 20250 14660 20256 14662
rect 19948 14651 20256 14660
rect 20608 14172 20916 14181
rect 20608 14170 20614 14172
rect 20670 14170 20694 14172
rect 20750 14170 20774 14172
rect 20830 14170 20854 14172
rect 20910 14170 20916 14172
rect 20670 14118 20672 14170
rect 20852 14118 20854 14170
rect 20608 14116 20614 14118
rect 20670 14116 20694 14118
rect 20750 14116 20774 14118
rect 20830 14116 20854 14118
rect 20910 14116 20916 14118
rect 20608 14107 20916 14116
rect 19948 13628 20256 13637
rect 19948 13626 19954 13628
rect 20010 13626 20034 13628
rect 20090 13626 20114 13628
rect 20170 13626 20194 13628
rect 20250 13626 20256 13628
rect 20010 13574 20012 13626
rect 20192 13574 20194 13626
rect 19948 13572 19954 13574
rect 20010 13572 20034 13574
rect 20090 13572 20114 13574
rect 20170 13572 20194 13574
rect 20250 13572 20256 13574
rect 19948 13563 20256 13572
rect 20608 13084 20916 13093
rect 20608 13082 20614 13084
rect 20670 13082 20694 13084
rect 20750 13082 20774 13084
rect 20830 13082 20854 13084
rect 20910 13082 20916 13084
rect 20670 13030 20672 13082
rect 20852 13030 20854 13082
rect 20608 13028 20614 13030
rect 20670 13028 20694 13030
rect 20750 13028 20774 13030
rect 20830 13028 20854 13030
rect 20910 13028 20916 13030
rect 20608 13019 20916 13028
rect 19948 12540 20256 12549
rect 19948 12538 19954 12540
rect 20010 12538 20034 12540
rect 20090 12538 20114 12540
rect 20170 12538 20194 12540
rect 20250 12538 20256 12540
rect 20010 12486 20012 12538
rect 20192 12486 20194 12538
rect 19948 12484 19954 12486
rect 20010 12484 20034 12486
rect 20090 12484 20114 12486
rect 20170 12484 20194 12486
rect 20250 12484 20256 12486
rect 19948 12475 20256 12484
rect 20608 11996 20916 12005
rect 20608 11994 20614 11996
rect 20670 11994 20694 11996
rect 20750 11994 20774 11996
rect 20830 11994 20854 11996
rect 20910 11994 20916 11996
rect 20670 11942 20672 11994
rect 20852 11942 20854 11994
rect 20608 11940 20614 11942
rect 20670 11940 20694 11942
rect 20750 11940 20774 11942
rect 20830 11940 20854 11942
rect 20910 11940 20916 11942
rect 20608 11931 20916 11940
rect 19948 11452 20256 11461
rect 19948 11450 19954 11452
rect 20010 11450 20034 11452
rect 20090 11450 20114 11452
rect 20170 11450 20194 11452
rect 20250 11450 20256 11452
rect 20010 11398 20012 11450
rect 20192 11398 20194 11450
rect 19948 11396 19954 11398
rect 20010 11396 20034 11398
rect 20090 11396 20114 11398
rect 20170 11396 20194 11398
rect 20250 11396 20256 11398
rect 19948 11387 20256 11396
rect 20608 10908 20916 10917
rect 20608 10906 20614 10908
rect 20670 10906 20694 10908
rect 20750 10906 20774 10908
rect 20830 10906 20854 10908
rect 20910 10906 20916 10908
rect 20670 10854 20672 10906
rect 20852 10854 20854 10906
rect 20608 10852 20614 10854
rect 20670 10852 20694 10854
rect 20750 10852 20774 10854
rect 20830 10852 20854 10854
rect 20910 10852 20916 10854
rect 20608 10843 20916 10852
rect 18880 10668 18932 10674
rect 18880 10610 18932 10616
rect 18892 10266 18920 10610
rect 22376 10464 22428 10470
rect 22376 10406 22428 10412
rect 19948 10364 20256 10373
rect 19948 10362 19954 10364
rect 20010 10362 20034 10364
rect 20090 10362 20114 10364
rect 20170 10362 20194 10364
rect 20250 10362 20256 10364
rect 20010 10310 20012 10362
rect 20192 10310 20194 10362
rect 19948 10308 19954 10310
rect 20010 10308 20034 10310
rect 20090 10308 20114 10310
rect 20170 10308 20194 10310
rect 20250 10308 20256 10310
rect 19948 10299 20256 10308
rect 22388 10305 22416 10406
rect 22374 10296 22430 10305
rect 18880 10260 18932 10266
rect 22374 10231 22430 10240
rect 18880 10202 18932 10208
rect 18236 10056 18288 10062
rect 18236 9998 18288 10004
rect 18248 5302 18276 9998
rect 20608 9820 20916 9829
rect 20608 9818 20614 9820
rect 20670 9818 20694 9820
rect 20750 9818 20774 9820
rect 20830 9818 20854 9820
rect 20910 9818 20916 9820
rect 20670 9766 20672 9818
rect 20852 9766 20854 9818
rect 20608 9764 20614 9766
rect 20670 9764 20694 9766
rect 20750 9764 20774 9766
rect 20830 9764 20854 9766
rect 20910 9764 20916 9766
rect 20608 9755 20916 9764
rect 19948 9276 20256 9285
rect 19948 9274 19954 9276
rect 20010 9274 20034 9276
rect 20090 9274 20114 9276
rect 20170 9274 20194 9276
rect 20250 9274 20256 9276
rect 20010 9222 20012 9274
rect 20192 9222 20194 9274
rect 19948 9220 19954 9222
rect 20010 9220 20034 9222
rect 20090 9220 20114 9222
rect 20170 9220 20194 9222
rect 20250 9220 20256 9222
rect 19948 9211 20256 9220
rect 20608 8732 20916 8741
rect 20608 8730 20614 8732
rect 20670 8730 20694 8732
rect 20750 8730 20774 8732
rect 20830 8730 20854 8732
rect 20910 8730 20916 8732
rect 20670 8678 20672 8730
rect 20852 8678 20854 8730
rect 20608 8676 20614 8678
rect 20670 8676 20694 8678
rect 20750 8676 20774 8678
rect 20830 8676 20854 8678
rect 20910 8676 20916 8678
rect 20608 8667 20916 8676
rect 19948 8188 20256 8197
rect 19948 8186 19954 8188
rect 20010 8186 20034 8188
rect 20090 8186 20114 8188
rect 20170 8186 20194 8188
rect 20250 8186 20256 8188
rect 20010 8134 20012 8186
rect 20192 8134 20194 8186
rect 19948 8132 19954 8134
rect 20010 8132 20034 8134
rect 20090 8132 20114 8134
rect 20170 8132 20194 8134
rect 20250 8132 20256 8134
rect 19948 8123 20256 8132
rect 20608 7644 20916 7653
rect 20608 7642 20614 7644
rect 20670 7642 20694 7644
rect 20750 7642 20774 7644
rect 20830 7642 20854 7644
rect 20910 7642 20916 7644
rect 20670 7590 20672 7642
rect 20852 7590 20854 7642
rect 20608 7588 20614 7590
rect 20670 7588 20694 7590
rect 20750 7588 20774 7590
rect 20830 7588 20854 7590
rect 20910 7588 20916 7590
rect 20608 7579 20916 7588
rect 19948 7100 20256 7109
rect 19948 7098 19954 7100
rect 20010 7098 20034 7100
rect 20090 7098 20114 7100
rect 20170 7098 20194 7100
rect 20250 7098 20256 7100
rect 20010 7046 20012 7098
rect 20192 7046 20194 7098
rect 19948 7044 19954 7046
rect 20010 7044 20034 7046
rect 20090 7044 20114 7046
rect 20170 7044 20194 7046
rect 20250 7044 20256 7046
rect 19948 7035 20256 7044
rect 20608 6556 20916 6565
rect 20608 6554 20614 6556
rect 20670 6554 20694 6556
rect 20750 6554 20774 6556
rect 20830 6554 20854 6556
rect 20910 6554 20916 6556
rect 20670 6502 20672 6554
rect 20852 6502 20854 6554
rect 20608 6500 20614 6502
rect 20670 6500 20694 6502
rect 20750 6500 20774 6502
rect 20830 6500 20854 6502
rect 20910 6500 20916 6502
rect 20608 6491 20916 6500
rect 19948 6012 20256 6021
rect 19948 6010 19954 6012
rect 20010 6010 20034 6012
rect 20090 6010 20114 6012
rect 20170 6010 20194 6012
rect 20250 6010 20256 6012
rect 20010 5958 20012 6010
rect 20192 5958 20194 6010
rect 19948 5956 19954 5958
rect 20010 5956 20034 5958
rect 20090 5956 20114 5958
rect 20170 5956 20194 5958
rect 20250 5956 20256 5958
rect 19948 5947 20256 5956
rect 20608 5468 20916 5477
rect 20608 5466 20614 5468
rect 20670 5466 20694 5468
rect 20750 5466 20774 5468
rect 20830 5466 20854 5468
rect 20910 5466 20916 5468
rect 20670 5414 20672 5466
rect 20852 5414 20854 5466
rect 20608 5412 20614 5414
rect 20670 5412 20694 5414
rect 20750 5412 20774 5414
rect 20830 5412 20854 5414
rect 20910 5412 20916 5414
rect 20608 5403 20916 5412
rect 18236 5296 18288 5302
rect 18236 5238 18288 5244
rect 19948 4924 20256 4933
rect 19948 4922 19954 4924
rect 20010 4922 20034 4924
rect 20090 4922 20114 4924
rect 20170 4922 20194 4924
rect 20250 4922 20256 4924
rect 20010 4870 20012 4922
rect 20192 4870 20194 4922
rect 19948 4868 19954 4870
rect 20010 4868 20034 4870
rect 20090 4868 20114 4870
rect 20170 4868 20194 4870
rect 20250 4868 20256 4870
rect 19948 4859 20256 4868
rect 20608 4380 20916 4389
rect 20608 4378 20614 4380
rect 20670 4378 20694 4380
rect 20750 4378 20774 4380
rect 20830 4378 20854 4380
rect 20910 4378 20916 4380
rect 20670 4326 20672 4378
rect 20852 4326 20854 4378
rect 20608 4324 20614 4326
rect 20670 4324 20694 4326
rect 20750 4324 20774 4326
rect 20830 4324 20854 4326
rect 20910 4324 20916 4326
rect 20608 4315 20916 4324
rect 18144 4208 18196 4214
rect 18144 4150 18196 4156
rect 22100 4140 22152 4146
rect 22100 4082 22152 4088
rect 19948 3836 20256 3845
rect 19948 3834 19954 3836
rect 20010 3834 20034 3836
rect 20090 3834 20114 3836
rect 20170 3834 20194 3836
rect 20250 3834 20256 3836
rect 20010 3782 20012 3834
rect 20192 3782 20194 3834
rect 19948 3780 19954 3782
rect 20010 3780 20034 3782
rect 20090 3780 20114 3782
rect 20170 3780 20194 3782
rect 20250 3780 20256 3782
rect 19948 3771 20256 3780
rect 20608 3292 20916 3301
rect 20608 3290 20614 3292
rect 20670 3290 20694 3292
rect 20750 3290 20774 3292
rect 20830 3290 20854 3292
rect 20910 3290 20916 3292
rect 20670 3238 20672 3290
rect 20852 3238 20854 3290
rect 20608 3236 20614 3238
rect 20670 3236 20694 3238
rect 20750 3236 20774 3238
rect 20830 3236 20854 3238
rect 20910 3236 20916 3238
rect 20608 3227 20916 3236
rect 19948 2748 20256 2757
rect 19948 2746 19954 2748
rect 20010 2746 20034 2748
rect 20090 2746 20114 2748
rect 20170 2746 20194 2748
rect 20250 2746 20256 2748
rect 20010 2694 20012 2746
rect 20192 2694 20194 2746
rect 19948 2692 19954 2694
rect 20010 2692 20034 2694
rect 20090 2692 20114 2694
rect 20170 2692 20194 2694
rect 20250 2692 20256 2694
rect 19948 2683 20256 2692
rect 22112 2650 22140 4082
rect 22100 2644 22152 2650
rect 22100 2586 22152 2592
rect 8484 2440 8536 2446
rect 8484 2382 8536 2388
rect 17132 2440 17184 2446
rect 17132 2382 17184 2388
rect 20 2372 72 2378
rect 20 2314 72 2320
rect 22836 2372 22888 2378
rect 22836 2314 22888 2320
rect 32 800 60 2314
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 4324 2204 4632 2213
rect 4324 2202 4330 2204
rect 4386 2202 4410 2204
rect 4466 2202 4490 2204
rect 4546 2202 4570 2204
rect 4626 2202 4632 2204
rect 4386 2150 4388 2202
rect 4568 2150 4570 2202
rect 4324 2148 4330 2150
rect 4386 2148 4410 2150
rect 4466 2148 4490 2150
rect 4546 2148 4570 2150
rect 4626 2148 4632 2150
rect 4324 2139 4632 2148
rect 8404 800 8432 2246
rect 9752 2204 10060 2213
rect 9752 2202 9758 2204
rect 9814 2202 9838 2204
rect 9894 2202 9918 2204
rect 9974 2202 9998 2204
rect 10054 2202 10060 2204
rect 9814 2150 9816 2202
rect 9996 2150 9998 2202
rect 9752 2148 9758 2150
rect 9814 2148 9838 2150
rect 9894 2148 9918 2150
rect 9974 2148 9998 2150
rect 10054 2148 10060 2150
rect 9752 2139 10060 2148
rect 15180 2204 15488 2213
rect 15180 2202 15186 2204
rect 15242 2202 15266 2204
rect 15322 2202 15346 2204
rect 15402 2202 15426 2204
rect 15482 2202 15488 2204
rect 15242 2150 15244 2202
rect 15424 2150 15426 2202
rect 15180 2148 15186 2150
rect 15242 2148 15266 2150
rect 15322 2148 15346 2150
rect 15402 2148 15426 2150
rect 15482 2148 15488 2150
rect 15180 2139 15488 2148
rect 16776 800 16804 2246
rect 20608 2204 20916 2213
rect 20608 2202 20614 2204
rect 20670 2202 20694 2204
rect 20750 2202 20774 2204
rect 20830 2202 20854 2204
rect 20910 2202 20916 2204
rect 20670 2150 20672 2202
rect 20852 2150 20854 2202
rect 20608 2148 20614 2150
rect 20670 2148 20694 2150
rect 20750 2148 20774 2150
rect 20830 2148 20854 2150
rect 20910 2148 20916 2150
rect 20608 2139 20916 2148
rect 22848 1465 22876 2314
rect 22834 1456 22890 1465
rect 22834 1391 22890 1400
rect 18 0 74 800
rect 8390 0 8446 800
rect 16762 0 16818 800
<< via2 >>
rect 4330 21786 4386 21788
rect 4410 21786 4466 21788
rect 4490 21786 4546 21788
rect 4570 21786 4626 21788
rect 4330 21734 4376 21786
rect 4376 21734 4386 21786
rect 4410 21734 4440 21786
rect 4440 21734 4452 21786
rect 4452 21734 4466 21786
rect 4490 21734 4504 21786
rect 4504 21734 4516 21786
rect 4516 21734 4546 21786
rect 4570 21734 4580 21786
rect 4580 21734 4626 21786
rect 4330 21732 4386 21734
rect 4410 21732 4466 21734
rect 4490 21732 4546 21734
rect 4570 21732 4626 21734
rect 9758 21786 9814 21788
rect 9838 21786 9894 21788
rect 9918 21786 9974 21788
rect 9998 21786 10054 21788
rect 9758 21734 9804 21786
rect 9804 21734 9814 21786
rect 9838 21734 9868 21786
rect 9868 21734 9880 21786
rect 9880 21734 9894 21786
rect 9918 21734 9932 21786
rect 9932 21734 9944 21786
rect 9944 21734 9974 21786
rect 9998 21734 10008 21786
rect 10008 21734 10054 21786
rect 9758 21732 9814 21734
rect 9838 21732 9894 21734
rect 9918 21732 9974 21734
rect 9998 21732 10054 21734
rect 15186 21786 15242 21788
rect 15266 21786 15322 21788
rect 15346 21786 15402 21788
rect 15426 21786 15482 21788
rect 15186 21734 15232 21786
rect 15232 21734 15242 21786
rect 15266 21734 15296 21786
rect 15296 21734 15308 21786
rect 15308 21734 15322 21786
rect 15346 21734 15360 21786
rect 15360 21734 15372 21786
rect 15372 21734 15402 21786
rect 15426 21734 15436 21786
rect 15436 21734 15482 21786
rect 15186 21732 15242 21734
rect 15266 21732 15322 21734
rect 15346 21732 15402 21734
rect 15426 21732 15482 21734
rect 20614 21786 20670 21788
rect 20694 21786 20750 21788
rect 20774 21786 20830 21788
rect 20854 21786 20910 21788
rect 20614 21734 20660 21786
rect 20660 21734 20670 21786
rect 20694 21734 20724 21786
rect 20724 21734 20736 21786
rect 20736 21734 20750 21786
rect 20774 21734 20788 21786
rect 20788 21734 20800 21786
rect 20800 21734 20830 21786
rect 20854 21734 20864 21786
rect 20864 21734 20910 21786
rect 20614 21732 20670 21734
rect 20694 21732 20750 21734
rect 20774 21732 20830 21734
rect 20854 21732 20910 21734
rect 3670 21242 3726 21244
rect 3750 21242 3806 21244
rect 3830 21242 3886 21244
rect 3910 21242 3966 21244
rect 3670 21190 3716 21242
rect 3716 21190 3726 21242
rect 3750 21190 3780 21242
rect 3780 21190 3792 21242
rect 3792 21190 3806 21242
rect 3830 21190 3844 21242
rect 3844 21190 3856 21242
rect 3856 21190 3886 21242
rect 3910 21190 3920 21242
rect 3920 21190 3966 21242
rect 3670 21188 3726 21190
rect 3750 21188 3806 21190
rect 3830 21188 3886 21190
rect 3910 21188 3966 21190
rect 3670 20154 3726 20156
rect 3750 20154 3806 20156
rect 3830 20154 3886 20156
rect 3910 20154 3966 20156
rect 3670 20102 3716 20154
rect 3716 20102 3726 20154
rect 3750 20102 3780 20154
rect 3780 20102 3792 20154
rect 3792 20102 3806 20154
rect 3830 20102 3844 20154
rect 3844 20102 3856 20154
rect 3856 20102 3886 20154
rect 3910 20102 3920 20154
rect 3920 20102 3966 20154
rect 3670 20100 3726 20102
rect 3750 20100 3806 20102
rect 3830 20100 3886 20102
rect 3910 20100 3966 20102
rect 3670 19066 3726 19068
rect 3750 19066 3806 19068
rect 3830 19066 3886 19068
rect 3910 19066 3966 19068
rect 3670 19014 3716 19066
rect 3716 19014 3726 19066
rect 3750 19014 3780 19066
rect 3780 19014 3792 19066
rect 3792 19014 3806 19066
rect 3830 19014 3844 19066
rect 3844 19014 3856 19066
rect 3856 19014 3886 19066
rect 3910 19014 3920 19066
rect 3920 19014 3966 19066
rect 3670 19012 3726 19014
rect 3750 19012 3806 19014
rect 3830 19012 3886 19014
rect 3910 19012 3966 19014
rect 9098 21242 9154 21244
rect 9178 21242 9234 21244
rect 9258 21242 9314 21244
rect 9338 21242 9394 21244
rect 9098 21190 9144 21242
rect 9144 21190 9154 21242
rect 9178 21190 9208 21242
rect 9208 21190 9220 21242
rect 9220 21190 9234 21242
rect 9258 21190 9272 21242
rect 9272 21190 9284 21242
rect 9284 21190 9314 21242
rect 9338 21190 9348 21242
rect 9348 21190 9394 21242
rect 9098 21188 9154 21190
rect 9178 21188 9234 21190
rect 9258 21188 9314 21190
rect 9338 21188 9394 21190
rect 4330 20698 4386 20700
rect 4410 20698 4466 20700
rect 4490 20698 4546 20700
rect 4570 20698 4626 20700
rect 4330 20646 4376 20698
rect 4376 20646 4386 20698
rect 4410 20646 4440 20698
rect 4440 20646 4452 20698
rect 4452 20646 4466 20698
rect 4490 20646 4504 20698
rect 4504 20646 4516 20698
rect 4516 20646 4546 20698
rect 4570 20646 4580 20698
rect 4580 20646 4626 20698
rect 4330 20644 4386 20646
rect 4410 20644 4466 20646
rect 4490 20644 4546 20646
rect 4570 20644 4626 20646
rect 9758 20698 9814 20700
rect 9838 20698 9894 20700
rect 9918 20698 9974 20700
rect 9998 20698 10054 20700
rect 9758 20646 9804 20698
rect 9804 20646 9814 20698
rect 9838 20646 9868 20698
rect 9868 20646 9880 20698
rect 9880 20646 9894 20698
rect 9918 20646 9932 20698
rect 9932 20646 9944 20698
rect 9944 20646 9974 20698
rect 9998 20646 10008 20698
rect 10008 20646 10054 20698
rect 9758 20644 9814 20646
rect 9838 20644 9894 20646
rect 9918 20644 9974 20646
rect 9998 20644 10054 20646
rect 9098 20154 9154 20156
rect 9178 20154 9234 20156
rect 9258 20154 9314 20156
rect 9338 20154 9394 20156
rect 9098 20102 9144 20154
rect 9144 20102 9154 20154
rect 9178 20102 9208 20154
rect 9208 20102 9220 20154
rect 9220 20102 9234 20154
rect 9258 20102 9272 20154
rect 9272 20102 9284 20154
rect 9284 20102 9314 20154
rect 9338 20102 9348 20154
rect 9348 20102 9394 20154
rect 9098 20100 9154 20102
rect 9178 20100 9234 20102
rect 9258 20100 9314 20102
rect 9338 20100 9394 20102
rect 4330 19610 4386 19612
rect 4410 19610 4466 19612
rect 4490 19610 4546 19612
rect 4570 19610 4626 19612
rect 4330 19558 4376 19610
rect 4376 19558 4386 19610
rect 4410 19558 4440 19610
rect 4440 19558 4452 19610
rect 4452 19558 4466 19610
rect 4490 19558 4504 19610
rect 4504 19558 4516 19610
rect 4516 19558 4546 19610
rect 4570 19558 4580 19610
rect 4580 19558 4626 19610
rect 4330 19556 4386 19558
rect 4410 19556 4466 19558
rect 4490 19556 4546 19558
rect 4570 19556 4626 19558
rect 9758 19610 9814 19612
rect 9838 19610 9894 19612
rect 9918 19610 9974 19612
rect 9998 19610 10054 19612
rect 9758 19558 9804 19610
rect 9804 19558 9814 19610
rect 9838 19558 9868 19610
rect 9868 19558 9880 19610
rect 9880 19558 9894 19610
rect 9918 19558 9932 19610
rect 9932 19558 9944 19610
rect 9944 19558 9974 19610
rect 9998 19558 10008 19610
rect 10008 19558 10054 19610
rect 9758 19556 9814 19558
rect 9838 19556 9894 19558
rect 9918 19556 9974 19558
rect 9998 19556 10054 19558
rect 9098 19066 9154 19068
rect 9178 19066 9234 19068
rect 9258 19066 9314 19068
rect 9338 19066 9394 19068
rect 9098 19014 9144 19066
rect 9144 19014 9154 19066
rect 9178 19014 9208 19066
rect 9208 19014 9220 19066
rect 9220 19014 9234 19066
rect 9258 19014 9272 19066
rect 9272 19014 9284 19066
rect 9284 19014 9314 19066
rect 9338 19014 9348 19066
rect 9348 19014 9394 19066
rect 9098 19012 9154 19014
rect 9178 19012 9234 19014
rect 9258 19012 9314 19014
rect 9338 19012 9394 19014
rect 14526 21242 14582 21244
rect 14606 21242 14662 21244
rect 14686 21242 14742 21244
rect 14766 21242 14822 21244
rect 14526 21190 14572 21242
rect 14572 21190 14582 21242
rect 14606 21190 14636 21242
rect 14636 21190 14648 21242
rect 14648 21190 14662 21242
rect 14686 21190 14700 21242
rect 14700 21190 14712 21242
rect 14712 21190 14742 21242
rect 14766 21190 14776 21242
rect 14776 21190 14822 21242
rect 14526 21188 14582 21190
rect 14606 21188 14662 21190
rect 14686 21188 14742 21190
rect 14766 21188 14822 21190
rect 15186 20698 15242 20700
rect 15266 20698 15322 20700
rect 15346 20698 15402 20700
rect 15426 20698 15482 20700
rect 15186 20646 15232 20698
rect 15232 20646 15242 20698
rect 15266 20646 15296 20698
rect 15296 20646 15308 20698
rect 15308 20646 15322 20698
rect 15346 20646 15360 20698
rect 15360 20646 15372 20698
rect 15372 20646 15402 20698
rect 15426 20646 15436 20698
rect 15436 20646 15482 20698
rect 15186 20644 15242 20646
rect 15266 20644 15322 20646
rect 15346 20644 15402 20646
rect 15426 20644 15482 20646
rect 14526 20154 14582 20156
rect 14606 20154 14662 20156
rect 14686 20154 14742 20156
rect 14766 20154 14822 20156
rect 14526 20102 14572 20154
rect 14572 20102 14582 20154
rect 14606 20102 14636 20154
rect 14636 20102 14648 20154
rect 14648 20102 14662 20154
rect 14686 20102 14700 20154
rect 14700 20102 14712 20154
rect 14712 20102 14742 20154
rect 14766 20102 14776 20154
rect 14776 20102 14822 20154
rect 14526 20100 14582 20102
rect 14606 20100 14662 20102
rect 14686 20100 14742 20102
rect 14766 20100 14822 20102
rect 15186 19610 15242 19612
rect 15266 19610 15322 19612
rect 15346 19610 15402 19612
rect 15426 19610 15482 19612
rect 15186 19558 15232 19610
rect 15232 19558 15242 19610
rect 15266 19558 15296 19610
rect 15296 19558 15308 19610
rect 15308 19558 15322 19610
rect 15346 19558 15360 19610
rect 15360 19558 15372 19610
rect 15372 19558 15402 19610
rect 15426 19558 15436 19610
rect 15436 19558 15482 19610
rect 15186 19556 15242 19558
rect 15266 19556 15322 19558
rect 15346 19556 15402 19558
rect 15426 19556 15482 19558
rect 14526 19066 14582 19068
rect 14606 19066 14662 19068
rect 14686 19066 14742 19068
rect 14766 19066 14822 19068
rect 14526 19014 14572 19066
rect 14572 19014 14582 19066
rect 14606 19014 14636 19066
rect 14636 19014 14648 19066
rect 14648 19014 14662 19066
rect 14686 19014 14700 19066
rect 14700 19014 14712 19066
rect 14712 19014 14742 19066
rect 14766 19014 14776 19066
rect 14776 19014 14822 19066
rect 14526 19012 14582 19014
rect 14606 19012 14662 19014
rect 14686 19012 14742 19014
rect 14766 19012 14822 19014
rect 4330 18522 4386 18524
rect 4410 18522 4466 18524
rect 4490 18522 4546 18524
rect 4570 18522 4626 18524
rect 4330 18470 4376 18522
rect 4376 18470 4386 18522
rect 4410 18470 4440 18522
rect 4440 18470 4452 18522
rect 4452 18470 4466 18522
rect 4490 18470 4504 18522
rect 4504 18470 4516 18522
rect 4516 18470 4546 18522
rect 4570 18470 4580 18522
rect 4580 18470 4626 18522
rect 4330 18468 4386 18470
rect 4410 18468 4466 18470
rect 4490 18468 4546 18470
rect 4570 18468 4626 18470
rect 9758 18522 9814 18524
rect 9838 18522 9894 18524
rect 9918 18522 9974 18524
rect 9998 18522 10054 18524
rect 9758 18470 9804 18522
rect 9804 18470 9814 18522
rect 9838 18470 9868 18522
rect 9868 18470 9880 18522
rect 9880 18470 9894 18522
rect 9918 18470 9932 18522
rect 9932 18470 9944 18522
rect 9944 18470 9974 18522
rect 9998 18470 10008 18522
rect 10008 18470 10054 18522
rect 9758 18468 9814 18470
rect 9838 18468 9894 18470
rect 9918 18468 9974 18470
rect 9998 18468 10054 18470
rect 15186 18522 15242 18524
rect 15266 18522 15322 18524
rect 15346 18522 15402 18524
rect 15426 18522 15482 18524
rect 15186 18470 15232 18522
rect 15232 18470 15242 18522
rect 15266 18470 15296 18522
rect 15296 18470 15308 18522
rect 15308 18470 15322 18522
rect 15346 18470 15360 18522
rect 15360 18470 15372 18522
rect 15372 18470 15402 18522
rect 15426 18470 15436 18522
rect 15436 18470 15482 18522
rect 15186 18468 15242 18470
rect 15266 18468 15322 18470
rect 15346 18468 15402 18470
rect 15426 18468 15482 18470
rect 3670 17978 3726 17980
rect 3750 17978 3806 17980
rect 3830 17978 3886 17980
rect 3910 17978 3966 17980
rect 3670 17926 3716 17978
rect 3716 17926 3726 17978
rect 3750 17926 3780 17978
rect 3780 17926 3792 17978
rect 3792 17926 3806 17978
rect 3830 17926 3844 17978
rect 3844 17926 3856 17978
rect 3856 17926 3886 17978
rect 3910 17926 3920 17978
rect 3920 17926 3966 17978
rect 3670 17924 3726 17926
rect 3750 17924 3806 17926
rect 3830 17924 3886 17926
rect 3910 17924 3966 17926
rect 1490 17856 1546 17912
rect 3670 16890 3726 16892
rect 3750 16890 3806 16892
rect 3830 16890 3886 16892
rect 3910 16890 3966 16892
rect 3670 16838 3716 16890
rect 3716 16838 3726 16890
rect 3750 16838 3780 16890
rect 3780 16838 3792 16890
rect 3792 16838 3806 16890
rect 3830 16838 3844 16890
rect 3844 16838 3856 16890
rect 3856 16838 3886 16890
rect 3910 16838 3920 16890
rect 3920 16838 3966 16890
rect 3670 16836 3726 16838
rect 3750 16836 3806 16838
rect 3830 16836 3886 16838
rect 3910 16836 3966 16838
rect 3670 15802 3726 15804
rect 3750 15802 3806 15804
rect 3830 15802 3886 15804
rect 3910 15802 3966 15804
rect 3670 15750 3716 15802
rect 3716 15750 3726 15802
rect 3750 15750 3780 15802
rect 3780 15750 3792 15802
rect 3792 15750 3806 15802
rect 3830 15750 3844 15802
rect 3844 15750 3856 15802
rect 3856 15750 3886 15802
rect 3910 15750 3920 15802
rect 3920 15750 3966 15802
rect 3670 15748 3726 15750
rect 3750 15748 3806 15750
rect 3830 15748 3886 15750
rect 3910 15748 3966 15750
rect 3670 14714 3726 14716
rect 3750 14714 3806 14716
rect 3830 14714 3886 14716
rect 3910 14714 3966 14716
rect 3670 14662 3716 14714
rect 3716 14662 3726 14714
rect 3750 14662 3780 14714
rect 3780 14662 3792 14714
rect 3792 14662 3806 14714
rect 3830 14662 3844 14714
rect 3844 14662 3856 14714
rect 3856 14662 3886 14714
rect 3910 14662 3920 14714
rect 3920 14662 3966 14714
rect 3670 14660 3726 14662
rect 3750 14660 3806 14662
rect 3830 14660 3886 14662
rect 3910 14660 3966 14662
rect 3670 13626 3726 13628
rect 3750 13626 3806 13628
rect 3830 13626 3886 13628
rect 3910 13626 3966 13628
rect 3670 13574 3716 13626
rect 3716 13574 3726 13626
rect 3750 13574 3780 13626
rect 3780 13574 3792 13626
rect 3792 13574 3806 13626
rect 3830 13574 3844 13626
rect 3844 13574 3856 13626
rect 3856 13574 3886 13626
rect 3910 13574 3920 13626
rect 3920 13574 3966 13626
rect 3670 13572 3726 13574
rect 3750 13572 3806 13574
rect 3830 13572 3886 13574
rect 3910 13572 3966 13574
rect 3670 12538 3726 12540
rect 3750 12538 3806 12540
rect 3830 12538 3886 12540
rect 3910 12538 3966 12540
rect 3670 12486 3716 12538
rect 3716 12486 3726 12538
rect 3750 12486 3780 12538
rect 3780 12486 3792 12538
rect 3792 12486 3806 12538
rect 3830 12486 3844 12538
rect 3844 12486 3856 12538
rect 3856 12486 3886 12538
rect 3910 12486 3920 12538
rect 3920 12486 3966 12538
rect 3670 12484 3726 12486
rect 3750 12484 3806 12486
rect 3830 12484 3886 12486
rect 3910 12484 3966 12486
rect 3670 11450 3726 11452
rect 3750 11450 3806 11452
rect 3830 11450 3886 11452
rect 3910 11450 3966 11452
rect 3670 11398 3716 11450
rect 3716 11398 3726 11450
rect 3750 11398 3780 11450
rect 3780 11398 3792 11450
rect 3792 11398 3806 11450
rect 3830 11398 3844 11450
rect 3844 11398 3856 11450
rect 3856 11398 3886 11450
rect 3910 11398 3920 11450
rect 3920 11398 3966 11450
rect 3670 11396 3726 11398
rect 3750 11396 3806 11398
rect 3830 11396 3886 11398
rect 3910 11396 3966 11398
rect 3670 10362 3726 10364
rect 3750 10362 3806 10364
rect 3830 10362 3886 10364
rect 3910 10362 3966 10364
rect 3670 10310 3716 10362
rect 3716 10310 3726 10362
rect 3750 10310 3780 10362
rect 3780 10310 3792 10362
rect 3792 10310 3806 10362
rect 3830 10310 3844 10362
rect 3844 10310 3856 10362
rect 3856 10310 3886 10362
rect 3910 10310 3920 10362
rect 3920 10310 3966 10362
rect 3670 10308 3726 10310
rect 3750 10308 3806 10310
rect 3830 10308 3886 10310
rect 3910 10308 3966 10310
rect 3670 9274 3726 9276
rect 3750 9274 3806 9276
rect 3830 9274 3886 9276
rect 3910 9274 3966 9276
rect 3670 9222 3716 9274
rect 3716 9222 3726 9274
rect 3750 9222 3780 9274
rect 3780 9222 3792 9274
rect 3792 9222 3806 9274
rect 3830 9222 3844 9274
rect 3844 9222 3856 9274
rect 3856 9222 3886 9274
rect 3910 9222 3920 9274
rect 3920 9222 3966 9274
rect 3670 9220 3726 9222
rect 3750 9220 3806 9222
rect 3830 9220 3886 9222
rect 3910 9220 3966 9222
rect 9098 17978 9154 17980
rect 9178 17978 9234 17980
rect 9258 17978 9314 17980
rect 9338 17978 9394 17980
rect 9098 17926 9144 17978
rect 9144 17926 9154 17978
rect 9178 17926 9208 17978
rect 9208 17926 9220 17978
rect 9220 17926 9234 17978
rect 9258 17926 9272 17978
rect 9272 17926 9284 17978
rect 9284 17926 9314 17978
rect 9338 17926 9348 17978
rect 9348 17926 9394 17978
rect 9098 17924 9154 17926
rect 9178 17924 9234 17926
rect 9258 17924 9314 17926
rect 9338 17924 9394 17926
rect 14526 17978 14582 17980
rect 14606 17978 14662 17980
rect 14686 17978 14742 17980
rect 14766 17978 14822 17980
rect 14526 17926 14572 17978
rect 14572 17926 14582 17978
rect 14606 17926 14636 17978
rect 14636 17926 14648 17978
rect 14648 17926 14662 17978
rect 14686 17926 14700 17978
rect 14700 17926 14712 17978
rect 14712 17926 14742 17978
rect 14766 17926 14776 17978
rect 14776 17926 14822 17978
rect 14526 17924 14582 17926
rect 14606 17924 14662 17926
rect 14686 17924 14742 17926
rect 14766 17924 14822 17926
rect 19954 21242 20010 21244
rect 20034 21242 20090 21244
rect 20114 21242 20170 21244
rect 20194 21242 20250 21244
rect 19954 21190 20000 21242
rect 20000 21190 20010 21242
rect 20034 21190 20064 21242
rect 20064 21190 20076 21242
rect 20076 21190 20090 21242
rect 20114 21190 20128 21242
rect 20128 21190 20140 21242
rect 20140 21190 20170 21242
rect 20194 21190 20204 21242
rect 20204 21190 20250 21242
rect 19954 21188 20010 21190
rect 20034 21188 20090 21190
rect 20114 21188 20170 21190
rect 20194 21188 20250 21190
rect 20614 20698 20670 20700
rect 20694 20698 20750 20700
rect 20774 20698 20830 20700
rect 20854 20698 20910 20700
rect 20614 20646 20660 20698
rect 20660 20646 20670 20698
rect 20694 20646 20724 20698
rect 20724 20646 20736 20698
rect 20736 20646 20750 20698
rect 20774 20646 20788 20698
rect 20788 20646 20800 20698
rect 20800 20646 20830 20698
rect 20854 20646 20864 20698
rect 20864 20646 20910 20698
rect 20614 20644 20670 20646
rect 20694 20644 20750 20646
rect 20774 20644 20830 20646
rect 20854 20644 20910 20646
rect 19954 20154 20010 20156
rect 20034 20154 20090 20156
rect 20114 20154 20170 20156
rect 20194 20154 20250 20156
rect 19954 20102 20000 20154
rect 20000 20102 20010 20154
rect 20034 20102 20064 20154
rect 20064 20102 20076 20154
rect 20076 20102 20090 20154
rect 20114 20102 20128 20154
rect 20128 20102 20140 20154
rect 20140 20102 20170 20154
rect 20194 20102 20204 20154
rect 20204 20102 20250 20154
rect 19954 20100 20010 20102
rect 20034 20100 20090 20102
rect 20114 20100 20170 20102
rect 20194 20100 20250 20102
rect 20614 19610 20670 19612
rect 20694 19610 20750 19612
rect 20774 19610 20830 19612
rect 20854 19610 20910 19612
rect 20614 19558 20660 19610
rect 20660 19558 20670 19610
rect 20694 19558 20724 19610
rect 20724 19558 20736 19610
rect 20736 19558 20750 19610
rect 20774 19558 20788 19610
rect 20788 19558 20800 19610
rect 20800 19558 20830 19610
rect 20854 19558 20864 19610
rect 20864 19558 20910 19610
rect 20614 19556 20670 19558
rect 20694 19556 20750 19558
rect 20774 19556 20830 19558
rect 20854 19556 20910 19558
rect 19954 19066 20010 19068
rect 20034 19066 20090 19068
rect 20114 19066 20170 19068
rect 20194 19066 20250 19068
rect 19954 19014 20000 19066
rect 20000 19014 20010 19066
rect 20034 19014 20064 19066
rect 20064 19014 20076 19066
rect 20076 19014 20090 19066
rect 20114 19014 20128 19066
rect 20128 19014 20140 19066
rect 20140 19014 20170 19066
rect 20194 19014 20204 19066
rect 20204 19014 20250 19066
rect 19954 19012 20010 19014
rect 20034 19012 20090 19014
rect 20114 19012 20170 19014
rect 20194 19012 20250 19014
rect 20614 18522 20670 18524
rect 20694 18522 20750 18524
rect 20774 18522 20830 18524
rect 20854 18522 20910 18524
rect 20614 18470 20660 18522
rect 20660 18470 20670 18522
rect 20694 18470 20724 18522
rect 20724 18470 20736 18522
rect 20736 18470 20750 18522
rect 20774 18470 20788 18522
rect 20788 18470 20800 18522
rect 20800 18470 20830 18522
rect 20854 18470 20864 18522
rect 20864 18470 20910 18522
rect 20614 18468 20670 18470
rect 20694 18468 20750 18470
rect 20774 18468 20830 18470
rect 20854 18468 20910 18470
rect 22834 19760 22890 19816
rect 19954 17978 20010 17980
rect 20034 17978 20090 17980
rect 20114 17978 20170 17980
rect 20194 17978 20250 17980
rect 19954 17926 20000 17978
rect 20000 17926 20010 17978
rect 20034 17926 20064 17978
rect 20064 17926 20076 17978
rect 20076 17926 20090 17978
rect 20114 17926 20128 17978
rect 20128 17926 20140 17978
rect 20140 17926 20170 17978
rect 20194 17926 20204 17978
rect 20204 17926 20250 17978
rect 19954 17924 20010 17926
rect 20034 17924 20090 17926
rect 20114 17924 20170 17926
rect 20194 17924 20250 17926
rect 4330 17434 4386 17436
rect 4410 17434 4466 17436
rect 4490 17434 4546 17436
rect 4570 17434 4626 17436
rect 4330 17382 4376 17434
rect 4376 17382 4386 17434
rect 4410 17382 4440 17434
rect 4440 17382 4452 17434
rect 4452 17382 4466 17434
rect 4490 17382 4504 17434
rect 4504 17382 4516 17434
rect 4516 17382 4546 17434
rect 4570 17382 4580 17434
rect 4580 17382 4626 17434
rect 4330 17380 4386 17382
rect 4410 17380 4466 17382
rect 4490 17380 4546 17382
rect 4570 17380 4626 17382
rect 9758 17434 9814 17436
rect 9838 17434 9894 17436
rect 9918 17434 9974 17436
rect 9998 17434 10054 17436
rect 9758 17382 9804 17434
rect 9804 17382 9814 17434
rect 9838 17382 9868 17434
rect 9868 17382 9880 17434
rect 9880 17382 9894 17434
rect 9918 17382 9932 17434
rect 9932 17382 9944 17434
rect 9944 17382 9974 17434
rect 9998 17382 10008 17434
rect 10008 17382 10054 17434
rect 9758 17380 9814 17382
rect 9838 17380 9894 17382
rect 9918 17380 9974 17382
rect 9998 17380 10054 17382
rect 15186 17434 15242 17436
rect 15266 17434 15322 17436
rect 15346 17434 15402 17436
rect 15426 17434 15482 17436
rect 15186 17382 15232 17434
rect 15232 17382 15242 17434
rect 15266 17382 15296 17434
rect 15296 17382 15308 17434
rect 15308 17382 15322 17434
rect 15346 17382 15360 17434
rect 15360 17382 15372 17434
rect 15372 17382 15402 17434
rect 15426 17382 15436 17434
rect 15436 17382 15482 17434
rect 15186 17380 15242 17382
rect 15266 17380 15322 17382
rect 15346 17380 15402 17382
rect 15426 17380 15482 17382
rect 9098 16890 9154 16892
rect 9178 16890 9234 16892
rect 9258 16890 9314 16892
rect 9338 16890 9394 16892
rect 9098 16838 9144 16890
rect 9144 16838 9154 16890
rect 9178 16838 9208 16890
rect 9208 16838 9220 16890
rect 9220 16838 9234 16890
rect 9258 16838 9272 16890
rect 9272 16838 9284 16890
rect 9284 16838 9314 16890
rect 9338 16838 9348 16890
rect 9348 16838 9394 16890
rect 9098 16836 9154 16838
rect 9178 16836 9234 16838
rect 9258 16836 9314 16838
rect 9338 16836 9394 16838
rect 14526 16890 14582 16892
rect 14606 16890 14662 16892
rect 14686 16890 14742 16892
rect 14766 16890 14822 16892
rect 14526 16838 14572 16890
rect 14572 16838 14582 16890
rect 14606 16838 14636 16890
rect 14636 16838 14648 16890
rect 14648 16838 14662 16890
rect 14686 16838 14700 16890
rect 14700 16838 14712 16890
rect 14712 16838 14742 16890
rect 14766 16838 14776 16890
rect 14776 16838 14822 16890
rect 14526 16836 14582 16838
rect 14606 16836 14662 16838
rect 14686 16836 14742 16838
rect 14766 16836 14822 16838
rect 4330 16346 4386 16348
rect 4410 16346 4466 16348
rect 4490 16346 4546 16348
rect 4570 16346 4626 16348
rect 4330 16294 4376 16346
rect 4376 16294 4386 16346
rect 4410 16294 4440 16346
rect 4440 16294 4452 16346
rect 4452 16294 4466 16346
rect 4490 16294 4504 16346
rect 4504 16294 4516 16346
rect 4516 16294 4546 16346
rect 4570 16294 4580 16346
rect 4580 16294 4626 16346
rect 4330 16292 4386 16294
rect 4410 16292 4466 16294
rect 4490 16292 4546 16294
rect 4570 16292 4626 16294
rect 9758 16346 9814 16348
rect 9838 16346 9894 16348
rect 9918 16346 9974 16348
rect 9998 16346 10054 16348
rect 9758 16294 9804 16346
rect 9804 16294 9814 16346
rect 9838 16294 9868 16346
rect 9868 16294 9880 16346
rect 9880 16294 9894 16346
rect 9918 16294 9932 16346
rect 9932 16294 9944 16346
rect 9944 16294 9974 16346
rect 9998 16294 10008 16346
rect 10008 16294 10054 16346
rect 9758 16292 9814 16294
rect 9838 16292 9894 16294
rect 9918 16292 9974 16294
rect 9998 16292 10054 16294
rect 15186 16346 15242 16348
rect 15266 16346 15322 16348
rect 15346 16346 15402 16348
rect 15426 16346 15482 16348
rect 15186 16294 15232 16346
rect 15232 16294 15242 16346
rect 15266 16294 15296 16346
rect 15296 16294 15308 16346
rect 15308 16294 15322 16346
rect 15346 16294 15360 16346
rect 15360 16294 15372 16346
rect 15372 16294 15402 16346
rect 15426 16294 15436 16346
rect 15436 16294 15482 16346
rect 15186 16292 15242 16294
rect 15266 16292 15322 16294
rect 15346 16292 15402 16294
rect 15426 16292 15482 16294
rect 9098 15802 9154 15804
rect 9178 15802 9234 15804
rect 9258 15802 9314 15804
rect 9338 15802 9394 15804
rect 9098 15750 9144 15802
rect 9144 15750 9154 15802
rect 9178 15750 9208 15802
rect 9208 15750 9220 15802
rect 9220 15750 9234 15802
rect 9258 15750 9272 15802
rect 9272 15750 9284 15802
rect 9284 15750 9314 15802
rect 9338 15750 9348 15802
rect 9348 15750 9394 15802
rect 9098 15748 9154 15750
rect 9178 15748 9234 15750
rect 9258 15748 9314 15750
rect 9338 15748 9394 15750
rect 14526 15802 14582 15804
rect 14606 15802 14662 15804
rect 14686 15802 14742 15804
rect 14766 15802 14822 15804
rect 14526 15750 14572 15802
rect 14572 15750 14582 15802
rect 14606 15750 14636 15802
rect 14636 15750 14648 15802
rect 14648 15750 14662 15802
rect 14686 15750 14700 15802
rect 14700 15750 14712 15802
rect 14712 15750 14742 15802
rect 14766 15750 14776 15802
rect 14776 15750 14822 15802
rect 14526 15748 14582 15750
rect 14606 15748 14662 15750
rect 14686 15748 14742 15750
rect 14766 15748 14822 15750
rect 4330 15258 4386 15260
rect 4410 15258 4466 15260
rect 4490 15258 4546 15260
rect 4570 15258 4626 15260
rect 4330 15206 4376 15258
rect 4376 15206 4386 15258
rect 4410 15206 4440 15258
rect 4440 15206 4452 15258
rect 4452 15206 4466 15258
rect 4490 15206 4504 15258
rect 4504 15206 4516 15258
rect 4516 15206 4546 15258
rect 4570 15206 4580 15258
rect 4580 15206 4626 15258
rect 4330 15204 4386 15206
rect 4410 15204 4466 15206
rect 4490 15204 4546 15206
rect 4570 15204 4626 15206
rect 9758 15258 9814 15260
rect 9838 15258 9894 15260
rect 9918 15258 9974 15260
rect 9998 15258 10054 15260
rect 9758 15206 9804 15258
rect 9804 15206 9814 15258
rect 9838 15206 9868 15258
rect 9868 15206 9880 15258
rect 9880 15206 9894 15258
rect 9918 15206 9932 15258
rect 9932 15206 9944 15258
rect 9944 15206 9974 15258
rect 9998 15206 10008 15258
rect 10008 15206 10054 15258
rect 9758 15204 9814 15206
rect 9838 15204 9894 15206
rect 9918 15204 9974 15206
rect 9998 15204 10054 15206
rect 15186 15258 15242 15260
rect 15266 15258 15322 15260
rect 15346 15258 15402 15260
rect 15426 15258 15482 15260
rect 15186 15206 15232 15258
rect 15232 15206 15242 15258
rect 15266 15206 15296 15258
rect 15296 15206 15308 15258
rect 15308 15206 15322 15258
rect 15346 15206 15360 15258
rect 15360 15206 15372 15258
rect 15372 15206 15402 15258
rect 15426 15206 15436 15258
rect 15436 15206 15482 15258
rect 15186 15204 15242 15206
rect 15266 15204 15322 15206
rect 15346 15204 15402 15206
rect 15426 15204 15482 15206
rect 9098 14714 9154 14716
rect 9178 14714 9234 14716
rect 9258 14714 9314 14716
rect 9338 14714 9394 14716
rect 9098 14662 9144 14714
rect 9144 14662 9154 14714
rect 9178 14662 9208 14714
rect 9208 14662 9220 14714
rect 9220 14662 9234 14714
rect 9258 14662 9272 14714
rect 9272 14662 9284 14714
rect 9284 14662 9314 14714
rect 9338 14662 9348 14714
rect 9348 14662 9394 14714
rect 9098 14660 9154 14662
rect 9178 14660 9234 14662
rect 9258 14660 9314 14662
rect 9338 14660 9394 14662
rect 14526 14714 14582 14716
rect 14606 14714 14662 14716
rect 14686 14714 14742 14716
rect 14766 14714 14822 14716
rect 14526 14662 14572 14714
rect 14572 14662 14582 14714
rect 14606 14662 14636 14714
rect 14636 14662 14648 14714
rect 14648 14662 14662 14714
rect 14686 14662 14700 14714
rect 14700 14662 14712 14714
rect 14712 14662 14742 14714
rect 14766 14662 14776 14714
rect 14776 14662 14822 14714
rect 14526 14660 14582 14662
rect 14606 14660 14662 14662
rect 14686 14660 14742 14662
rect 14766 14660 14822 14662
rect 4330 14170 4386 14172
rect 4410 14170 4466 14172
rect 4490 14170 4546 14172
rect 4570 14170 4626 14172
rect 4330 14118 4376 14170
rect 4376 14118 4386 14170
rect 4410 14118 4440 14170
rect 4440 14118 4452 14170
rect 4452 14118 4466 14170
rect 4490 14118 4504 14170
rect 4504 14118 4516 14170
rect 4516 14118 4546 14170
rect 4570 14118 4580 14170
rect 4580 14118 4626 14170
rect 4330 14116 4386 14118
rect 4410 14116 4466 14118
rect 4490 14116 4546 14118
rect 4570 14116 4626 14118
rect 9758 14170 9814 14172
rect 9838 14170 9894 14172
rect 9918 14170 9974 14172
rect 9998 14170 10054 14172
rect 9758 14118 9804 14170
rect 9804 14118 9814 14170
rect 9838 14118 9868 14170
rect 9868 14118 9880 14170
rect 9880 14118 9894 14170
rect 9918 14118 9932 14170
rect 9932 14118 9944 14170
rect 9944 14118 9974 14170
rect 9998 14118 10008 14170
rect 10008 14118 10054 14170
rect 9758 14116 9814 14118
rect 9838 14116 9894 14118
rect 9918 14116 9974 14118
rect 9998 14116 10054 14118
rect 15186 14170 15242 14172
rect 15266 14170 15322 14172
rect 15346 14170 15402 14172
rect 15426 14170 15482 14172
rect 15186 14118 15232 14170
rect 15232 14118 15242 14170
rect 15266 14118 15296 14170
rect 15296 14118 15308 14170
rect 15308 14118 15322 14170
rect 15346 14118 15360 14170
rect 15360 14118 15372 14170
rect 15372 14118 15402 14170
rect 15426 14118 15436 14170
rect 15436 14118 15482 14170
rect 15186 14116 15242 14118
rect 15266 14116 15322 14118
rect 15346 14116 15402 14118
rect 15426 14116 15482 14118
rect 9098 13626 9154 13628
rect 9178 13626 9234 13628
rect 9258 13626 9314 13628
rect 9338 13626 9394 13628
rect 9098 13574 9144 13626
rect 9144 13574 9154 13626
rect 9178 13574 9208 13626
rect 9208 13574 9220 13626
rect 9220 13574 9234 13626
rect 9258 13574 9272 13626
rect 9272 13574 9284 13626
rect 9284 13574 9314 13626
rect 9338 13574 9348 13626
rect 9348 13574 9394 13626
rect 9098 13572 9154 13574
rect 9178 13572 9234 13574
rect 9258 13572 9314 13574
rect 9338 13572 9394 13574
rect 14526 13626 14582 13628
rect 14606 13626 14662 13628
rect 14686 13626 14742 13628
rect 14766 13626 14822 13628
rect 14526 13574 14572 13626
rect 14572 13574 14582 13626
rect 14606 13574 14636 13626
rect 14636 13574 14648 13626
rect 14648 13574 14662 13626
rect 14686 13574 14700 13626
rect 14700 13574 14712 13626
rect 14712 13574 14742 13626
rect 14766 13574 14776 13626
rect 14776 13574 14822 13626
rect 14526 13572 14582 13574
rect 14606 13572 14662 13574
rect 14686 13572 14742 13574
rect 14766 13572 14822 13574
rect 4330 13082 4386 13084
rect 4410 13082 4466 13084
rect 4490 13082 4546 13084
rect 4570 13082 4626 13084
rect 4330 13030 4376 13082
rect 4376 13030 4386 13082
rect 4410 13030 4440 13082
rect 4440 13030 4452 13082
rect 4452 13030 4466 13082
rect 4490 13030 4504 13082
rect 4504 13030 4516 13082
rect 4516 13030 4546 13082
rect 4570 13030 4580 13082
rect 4580 13030 4626 13082
rect 4330 13028 4386 13030
rect 4410 13028 4466 13030
rect 4490 13028 4546 13030
rect 4570 13028 4626 13030
rect 9758 13082 9814 13084
rect 9838 13082 9894 13084
rect 9918 13082 9974 13084
rect 9998 13082 10054 13084
rect 9758 13030 9804 13082
rect 9804 13030 9814 13082
rect 9838 13030 9868 13082
rect 9868 13030 9880 13082
rect 9880 13030 9894 13082
rect 9918 13030 9932 13082
rect 9932 13030 9944 13082
rect 9944 13030 9974 13082
rect 9998 13030 10008 13082
rect 10008 13030 10054 13082
rect 9758 13028 9814 13030
rect 9838 13028 9894 13030
rect 9918 13028 9974 13030
rect 9998 13028 10054 13030
rect 15186 13082 15242 13084
rect 15266 13082 15322 13084
rect 15346 13082 15402 13084
rect 15426 13082 15482 13084
rect 15186 13030 15232 13082
rect 15232 13030 15242 13082
rect 15266 13030 15296 13082
rect 15296 13030 15308 13082
rect 15308 13030 15322 13082
rect 15346 13030 15360 13082
rect 15360 13030 15372 13082
rect 15372 13030 15402 13082
rect 15426 13030 15436 13082
rect 15436 13030 15482 13082
rect 15186 13028 15242 13030
rect 15266 13028 15322 13030
rect 15346 13028 15402 13030
rect 15426 13028 15482 13030
rect 9098 12538 9154 12540
rect 9178 12538 9234 12540
rect 9258 12538 9314 12540
rect 9338 12538 9394 12540
rect 9098 12486 9144 12538
rect 9144 12486 9154 12538
rect 9178 12486 9208 12538
rect 9208 12486 9220 12538
rect 9220 12486 9234 12538
rect 9258 12486 9272 12538
rect 9272 12486 9284 12538
rect 9284 12486 9314 12538
rect 9338 12486 9348 12538
rect 9348 12486 9394 12538
rect 9098 12484 9154 12486
rect 9178 12484 9234 12486
rect 9258 12484 9314 12486
rect 9338 12484 9394 12486
rect 14526 12538 14582 12540
rect 14606 12538 14662 12540
rect 14686 12538 14742 12540
rect 14766 12538 14822 12540
rect 14526 12486 14572 12538
rect 14572 12486 14582 12538
rect 14606 12486 14636 12538
rect 14636 12486 14648 12538
rect 14648 12486 14662 12538
rect 14686 12486 14700 12538
rect 14700 12486 14712 12538
rect 14712 12486 14742 12538
rect 14766 12486 14776 12538
rect 14776 12486 14822 12538
rect 14526 12484 14582 12486
rect 14606 12484 14662 12486
rect 14686 12484 14742 12486
rect 14766 12484 14822 12486
rect 4330 11994 4386 11996
rect 4410 11994 4466 11996
rect 4490 11994 4546 11996
rect 4570 11994 4626 11996
rect 4330 11942 4376 11994
rect 4376 11942 4386 11994
rect 4410 11942 4440 11994
rect 4440 11942 4452 11994
rect 4452 11942 4466 11994
rect 4490 11942 4504 11994
rect 4504 11942 4516 11994
rect 4516 11942 4546 11994
rect 4570 11942 4580 11994
rect 4580 11942 4626 11994
rect 4330 11940 4386 11942
rect 4410 11940 4466 11942
rect 4490 11940 4546 11942
rect 4570 11940 4626 11942
rect 9758 11994 9814 11996
rect 9838 11994 9894 11996
rect 9918 11994 9974 11996
rect 9998 11994 10054 11996
rect 9758 11942 9804 11994
rect 9804 11942 9814 11994
rect 9838 11942 9868 11994
rect 9868 11942 9880 11994
rect 9880 11942 9894 11994
rect 9918 11942 9932 11994
rect 9932 11942 9944 11994
rect 9944 11942 9974 11994
rect 9998 11942 10008 11994
rect 10008 11942 10054 11994
rect 9758 11940 9814 11942
rect 9838 11940 9894 11942
rect 9918 11940 9974 11942
rect 9998 11940 10054 11942
rect 15186 11994 15242 11996
rect 15266 11994 15322 11996
rect 15346 11994 15402 11996
rect 15426 11994 15482 11996
rect 15186 11942 15232 11994
rect 15232 11942 15242 11994
rect 15266 11942 15296 11994
rect 15296 11942 15308 11994
rect 15308 11942 15322 11994
rect 15346 11942 15360 11994
rect 15360 11942 15372 11994
rect 15372 11942 15402 11994
rect 15426 11942 15436 11994
rect 15436 11942 15482 11994
rect 15186 11940 15242 11942
rect 15266 11940 15322 11942
rect 15346 11940 15402 11942
rect 15426 11940 15482 11942
rect 9098 11450 9154 11452
rect 9178 11450 9234 11452
rect 9258 11450 9314 11452
rect 9338 11450 9394 11452
rect 9098 11398 9144 11450
rect 9144 11398 9154 11450
rect 9178 11398 9208 11450
rect 9208 11398 9220 11450
rect 9220 11398 9234 11450
rect 9258 11398 9272 11450
rect 9272 11398 9284 11450
rect 9284 11398 9314 11450
rect 9338 11398 9348 11450
rect 9348 11398 9394 11450
rect 9098 11396 9154 11398
rect 9178 11396 9234 11398
rect 9258 11396 9314 11398
rect 9338 11396 9394 11398
rect 14526 11450 14582 11452
rect 14606 11450 14662 11452
rect 14686 11450 14742 11452
rect 14766 11450 14822 11452
rect 14526 11398 14572 11450
rect 14572 11398 14582 11450
rect 14606 11398 14636 11450
rect 14636 11398 14648 11450
rect 14648 11398 14662 11450
rect 14686 11398 14700 11450
rect 14700 11398 14712 11450
rect 14712 11398 14742 11450
rect 14766 11398 14776 11450
rect 14776 11398 14822 11450
rect 14526 11396 14582 11398
rect 14606 11396 14662 11398
rect 14686 11396 14742 11398
rect 14766 11396 14822 11398
rect 4330 10906 4386 10908
rect 4410 10906 4466 10908
rect 4490 10906 4546 10908
rect 4570 10906 4626 10908
rect 4330 10854 4376 10906
rect 4376 10854 4386 10906
rect 4410 10854 4440 10906
rect 4440 10854 4452 10906
rect 4452 10854 4466 10906
rect 4490 10854 4504 10906
rect 4504 10854 4516 10906
rect 4516 10854 4546 10906
rect 4570 10854 4580 10906
rect 4580 10854 4626 10906
rect 4330 10852 4386 10854
rect 4410 10852 4466 10854
rect 4490 10852 4546 10854
rect 4570 10852 4626 10854
rect 9758 10906 9814 10908
rect 9838 10906 9894 10908
rect 9918 10906 9974 10908
rect 9998 10906 10054 10908
rect 9758 10854 9804 10906
rect 9804 10854 9814 10906
rect 9838 10854 9868 10906
rect 9868 10854 9880 10906
rect 9880 10854 9894 10906
rect 9918 10854 9932 10906
rect 9932 10854 9944 10906
rect 9944 10854 9974 10906
rect 9998 10854 10008 10906
rect 10008 10854 10054 10906
rect 9758 10852 9814 10854
rect 9838 10852 9894 10854
rect 9918 10852 9974 10854
rect 9998 10852 10054 10854
rect 15186 10906 15242 10908
rect 15266 10906 15322 10908
rect 15346 10906 15402 10908
rect 15426 10906 15482 10908
rect 15186 10854 15232 10906
rect 15232 10854 15242 10906
rect 15266 10854 15296 10906
rect 15296 10854 15308 10906
rect 15308 10854 15322 10906
rect 15346 10854 15360 10906
rect 15360 10854 15372 10906
rect 15372 10854 15402 10906
rect 15426 10854 15436 10906
rect 15436 10854 15482 10906
rect 15186 10852 15242 10854
rect 15266 10852 15322 10854
rect 15346 10852 15402 10854
rect 15426 10852 15482 10854
rect 9098 10362 9154 10364
rect 9178 10362 9234 10364
rect 9258 10362 9314 10364
rect 9338 10362 9394 10364
rect 9098 10310 9144 10362
rect 9144 10310 9154 10362
rect 9178 10310 9208 10362
rect 9208 10310 9220 10362
rect 9220 10310 9234 10362
rect 9258 10310 9272 10362
rect 9272 10310 9284 10362
rect 9284 10310 9314 10362
rect 9338 10310 9348 10362
rect 9348 10310 9394 10362
rect 9098 10308 9154 10310
rect 9178 10308 9234 10310
rect 9258 10308 9314 10310
rect 9338 10308 9394 10310
rect 14526 10362 14582 10364
rect 14606 10362 14662 10364
rect 14686 10362 14742 10364
rect 14766 10362 14822 10364
rect 14526 10310 14572 10362
rect 14572 10310 14582 10362
rect 14606 10310 14636 10362
rect 14636 10310 14648 10362
rect 14648 10310 14662 10362
rect 14686 10310 14700 10362
rect 14700 10310 14712 10362
rect 14712 10310 14742 10362
rect 14766 10310 14776 10362
rect 14776 10310 14822 10362
rect 14526 10308 14582 10310
rect 14606 10308 14662 10310
rect 14686 10308 14742 10310
rect 14766 10308 14822 10310
rect 4330 9818 4386 9820
rect 4410 9818 4466 9820
rect 4490 9818 4546 9820
rect 4570 9818 4626 9820
rect 4330 9766 4376 9818
rect 4376 9766 4386 9818
rect 4410 9766 4440 9818
rect 4440 9766 4452 9818
rect 4452 9766 4466 9818
rect 4490 9766 4504 9818
rect 4504 9766 4516 9818
rect 4516 9766 4546 9818
rect 4570 9766 4580 9818
rect 4580 9766 4626 9818
rect 4330 9764 4386 9766
rect 4410 9764 4466 9766
rect 4490 9764 4546 9766
rect 4570 9764 4626 9766
rect 9758 9818 9814 9820
rect 9838 9818 9894 9820
rect 9918 9818 9974 9820
rect 9998 9818 10054 9820
rect 9758 9766 9804 9818
rect 9804 9766 9814 9818
rect 9838 9766 9868 9818
rect 9868 9766 9880 9818
rect 9880 9766 9894 9818
rect 9918 9766 9932 9818
rect 9932 9766 9944 9818
rect 9944 9766 9974 9818
rect 9998 9766 10008 9818
rect 10008 9766 10054 9818
rect 9758 9764 9814 9766
rect 9838 9764 9894 9766
rect 9918 9764 9974 9766
rect 9998 9764 10054 9766
rect 15186 9818 15242 9820
rect 15266 9818 15322 9820
rect 15346 9818 15402 9820
rect 15426 9818 15482 9820
rect 15186 9766 15232 9818
rect 15232 9766 15242 9818
rect 15266 9766 15296 9818
rect 15296 9766 15308 9818
rect 15308 9766 15322 9818
rect 15346 9766 15360 9818
rect 15360 9766 15372 9818
rect 15372 9766 15402 9818
rect 15426 9766 15436 9818
rect 15436 9766 15482 9818
rect 15186 9764 15242 9766
rect 15266 9764 15322 9766
rect 15346 9764 15402 9766
rect 15426 9764 15482 9766
rect 9098 9274 9154 9276
rect 9178 9274 9234 9276
rect 9258 9274 9314 9276
rect 9338 9274 9394 9276
rect 9098 9222 9144 9274
rect 9144 9222 9154 9274
rect 9178 9222 9208 9274
rect 9208 9222 9220 9274
rect 9220 9222 9234 9274
rect 9258 9222 9272 9274
rect 9272 9222 9284 9274
rect 9284 9222 9314 9274
rect 9338 9222 9348 9274
rect 9348 9222 9394 9274
rect 9098 9220 9154 9222
rect 9178 9220 9234 9222
rect 9258 9220 9314 9222
rect 9338 9220 9394 9222
rect 14526 9274 14582 9276
rect 14606 9274 14662 9276
rect 14686 9274 14742 9276
rect 14766 9274 14822 9276
rect 14526 9222 14572 9274
rect 14572 9222 14582 9274
rect 14606 9222 14636 9274
rect 14636 9222 14648 9274
rect 14648 9222 14662 9274
rect 14686 9222 14700 9274
rect 14700 9222 14712 9274
rect 14712 9222 14742 9274
rect 14766 9222 14776 9274
rect 14776 9222 14822 9274
rect 14526 9220 14582 9222
rect 14606 9220 14662 9222
rect 14686 9220 14742 9222
rect 14766 9220 14822 9222
rect 938 8900 994 8936
rect 938 8880 940 8900
rect 940 8880 992 8900
rect 992 8880 994 8900
rect 3670 8186 3726 8188
rect 3750 8186 3806 8188
rect 3830 8186 3886 8188
rect 3910 8186 3966 8188
rect 3670 8134 3716 8186
rect 3716 8134 3726 8186
rect 3750 8134 3780 8186
rect 3780 8134 3792 8186
rect 3792 8134 3806 8186
rect 3830 8134 3844 8186
rect 3844 8134 3856 8186
rect 3856 8134 3886 8186
rect 3910 8134 3920 8186
rect 3920 8134 3966 8186
rect 3670 8132 3726 8134
rect 3750 8132 3806 8134
rect 3830 8132 3886 8134
rect 3910 8132 3966 8134
rect 3670 7098 3726 7100
rect 3750 7098 3806 7100
rect 3830 7098 3886 7100
rect 3910 7098 3966 7100
rect 3670 7046 3716 7098
rect 3716 7046 3726 7098
rect 3750 7046 3780 7098
rect 3780 7046 3792 7098
rect 3792 7046 3806 7098
rect 3830 7046 3844 7098
rect 3844 7046 3856 7098
rect 3856 7046 3886 7098
rect 3910 7046 3920 7098
rect 3920 7046 3966 7098
rect 3670 7044 3726 7046
rect 3750 7044 3806 7046
rect 3830 7044 3886 7046
rect 3910 7044 3966 7046
rect 3670 6010 3726 6012
rect 3750 6010 3806 6012
rect 3830 6010 3886 6012
rect 3910 6010 3966 6012
rect 3670 5958 3716 6010
rect 3716 5958 3726 6010
rect 3750 5958 3780 6010
rect 3780 5958 3792 6010
rect 3792 5958 3806 6010
rect 3830 5958 3844 6010
rect 3844 5958 3856 6010
rect 3856 5958 3886 6010
rect 3910 5958 3920 6010
rect 3920 5958 3966 6010
rect 3670 5956 3726 5958
rect 3750 5956 3806 5958
rect 3830 5956 3886 5958
rect 3910 5956 3966 5958
rect 3670 4922 3726 4924
rect 3750 4922 3806 4924
rect 3830 4922 3886 4924
rect 3910 4922 3966 4924
rect 3670 4870 3716 4922
rect 3716 4870 3726 4922
rect 3750 4870 3780 4922
rect 3780 4870 3792 4922
rect 3792 4870 3806 4922
rect 3830 4870 3844 4922
rect 3844 4870 3856 4922
rect 3856 4870 3886 4922
rect 3910 4870 3920 4922
rect 3920 4870 3966 4922
rect 3670 4868 3726 4870
rect 3750 4868 3806 4870
rect 3830 4868 3886 4870
rect 3910 4868 3966 4870
rect 4330 8730 4386 8732
rect 4410 8730 4466 8732
rect 4490 8730 4546 8732
rect 4570 8730 4626 8732
rect 4330 8678 4376 8730
rect 4376 8678 4386 8730
rect 4410 8678 4440 8730
rect 4440 8678 4452 8730
rect 4452 8678 4466 8730
rect 4490 8678 4504 8730
rect 4504 8678 4516 8730
rect 4516 8678 4546 8730
rect 4570 8678 4580 8730
rect 4580 8678 4626 8730
rect 4330 8676 4386 8678
rect 4410 8676 4466 8678
rect 4490 8676 4546 8678
rect 4570 8676 4626 8678
rect 4330 7642 4386 7644
rect 4410 7642 4466 7644
rect 4490 7642 4546 7644
rect 4570 7642 4626 7644
rect 4330 7590 4376 7642
rect 4376 7590 4386 7642
rect 4410 7590 4440 7642
rect 4440 7590 4452 7642
rect 4452 7590 4466 7642
rect 4490 7590 4504 7642
rect 4504 7590 4516 7642
rect 4516 7590 4546 7642
rect 4570 7590 4580 7642
rect 4580 7590 4626 7642
rect 4330 7588 4386 7590
rect 4410 7588 4466 7590
rect 4490 7588 4546 7590
rect 4570 7588 4626 7590
rect 4330 6554 4386 6556
rect 4410 6554 4466 6556
rect 4490 6554 4546 6556
rect 4570 6554 4626 6556
rect 4330 6502 4376 6554
rect 4376 6502 4386 6554
rect 4410 6502 4440 6554
rect 4440 6502 4452 6554
rect 4452 6502 4466 6554
rect 4490 6502 4504 6554
rect 4504 6502 4516 6554
rect 4516 6502 4546 6554
rect 4570 6502 4580 6554
rect 4580 6502 4626 6554
rect 4330 6500 4386 6502
rect 4410 6500 4466 6502
rect 4490 6500 4546 6502
rect 4570 6500 4626 6502
rect 4330 5466 4386 5468
rect 4410 5466 4466 5468
rect 4490 5466 4546 5468
rect 4570 5466 4626 5468
rect 4330 5414 4376 5466
rect 4376 5414 4386 5466
rect 4410 5414 4440 5466
rect 4440 5414 4452 5466
rect 4452 5414 4466 5466
rect 4490 5414 4504 5466
rect 4504 5414 4516 5466
rect 4516 5414 4546 5466
rect 4570 5414 4580 5466
rect 4580 5414 4626 5466
rect 4330 5412 4386 5414
rect 4410 5412 4466 5414
rect 4490 5412 4546 5414
rect 4570 5412 4626 5414
rect 4330 4378 4386 4380
rect 4410 4378 4466 4380
rect 4490 4378 4546 4380
rect 4570 4378 4626 4380
rect 4330 4326 4376 4378
rect 4376 4326 4386 4378
rect 4410 4326 4440 4378
rect 4440 4326 4452 4378
rect 4452 4326 4466 4378
rect 4490 4326 4504 4378
rect 4504 4326 4516 4378
rect 4516 4326 4546 4378
rect 4570 4326 4580 4378
rect 4580 4326 4626 4378
rect 4330 4324 4386 4326
rect 4410 4324 4466 4326
rect 4490 4324 4546 4326
rect 4570 4324 4626 4326
rect 9758 8730 9814 8732
rect 9838 8730 9894 8732
rect 9918 8730 9974 8732
rect 9998 8730 10054 8732
rect 9758 8678 9804 8730
rect 9804 8678 9814 8730
rect 9838 8678 9868 8730
rect 9868 8678 9880 8730
rect 9880 8678 9894 8730
rect 9918 8678 9932 8730
rect 9932 8678 9944 8730
rect 9944 8678 9974 8730
rect 9998 8678 10008 8730
rect 10008 8678 10054 8730
rect 9758 8676 9814 8678
rect 9838 8676 9894 8678
rect 9918 8676 9974 8678
rect 9998 8676 10054 8678
rect 15186 8730 15242 8732
rect 15266 8730 15322 8732
rect 15346 8730 15402 8732
rect 15426 8730 15482 8732
rect 15186 8678 15232 8730
rect 15232 8678 15242 8730
rect 15266 8678 15296 8730
rect 15296 8678 15308 8730
rect 15308 8678 15322 8730
rect 15346 8678 15360 8730
rect 15360 8678 15372 8730
rect 15372 8678 15402 8730
rect 15426 8678 15436 8730
rect 15436 8678 15482 8730
rect 15186 8676 15242 8678
rect 15266 8676 15322 8678
rect 15346 8676 15402 8678
rect 15426 8676 15482 8678
rect 9098 8186 9154 8188
rect 9178 8186 9234 8188
rect 9258 8186 9314 8188
rect 9338 8186 9394 8188
rect 9098 8134 9144 8186
rect 9144 8134 9154 8186
rect 9178 8134 9208 8186
rect 9208 8134 9220 8186
rect 9220 8134 9234 8186
rect 9258 8134 9272 8186
rect 9272 8134 9284 8186
rect 9284 8134 9314 8186
rect 9338 8134 9348 8186
rect 9348 8134 9394 8186
rect 9098 8132 9154 8134
rect 9178 8132 9234 8134
rect 9258 8132 9314 8134
rect 9338 8132 9394 8134
rect 14526 8186 14582 8188
rect 14606 8186 14662 8188
rect 14686 8186 14742 8188
rect 14766 8186 14822 8188
rect 14526 8134 14572 8186
rect 14572 8134 14582 8186
rect 14606 8134 14636 8186
rect 14636 8134 14648 8186
rect 14648 8134 14662 8186
rect 14686 8134 14700 8186
rect 14700 8134 14712 8186
rect 14712 8134 14742 8186
rect 14766 8134 14776 8186
rect 14776 8134 14822 8186
rect 14526 8132 14582 8134
rect 14606 8132 14662 8134
rect 14686 8132 14742 8134
rect 14766 8132 14822 8134
rect 9758 7642 9814 7644
rect 9838 7642 9894 7644
rect 9918 7642 9974 7644
rect 9998 7642 10054 7644
rect 9758 7590 9804 7642
rect 9804 7590 9814 7642
rect 9838 7590 9868 7642
rect 9868 7590 9880 7642
rect 9880 7590 9894 7642
rect 9918 7590 9932 7642
rect 9932 7590 9944 7642
rect 9944 7590 9974 7642
rect 9998 7590 10008 7642
rect 10008 7590 10054 7642
rect 9758 7588 9814 7590
rect 9838 7588 9894 7590
rect 9918 7588 9974 7590
rect 9998 7588 10054 7590
rect 15186 7642 15242 7644
rect 15266 7642 15322 7644
rect 15346 7642 15402 7644
rect 15426 7642 15482 7644
rect 15186 7590 15232 7642
rect 15232 7590 15242 7642
rect 15266 7590 15296 7642
rect 15296 7590 15308 7642
rect 15308 7590 15322 7642
rect 15346 7590 15360 7642
rect 15360 7590 15372 7642
rect 15372 7590 15402 7642
rect 15426 7590 15436 7642
rect 15436 7590 15482 7642
rect 15186 7588 15242 7590
rect 15266 7588 15322 7590
rect 15346 7588 15402 7590
rect 15426 7588 15482 7590
rect 9098 7098 9154 7100
rect 9178 7098 9234 7100
rect 9258 7098 9314 7100
rect 9338 7098 9394 7100
rect 9098 7046 9144 7098
rect 9144 7046 9154 7098
rect 9178 7046 9208 7098
rect 9208 7046 9220 7098
rect 9220 7046 9234 7098
rect 9258 7046 9272 7098
rect 9272 7046 9284 7098
rect 9284 7046 9314 7098
rect 9338 7046 9348 7098
rect 9348 7046 9394 7098
rect 9098 7044 9154 7046
rect 9178 7044 9234 7046
rect 9258 7044 9314 7046
rect 9338 7044 9394 7046
rect 14526 7098 14582 7100
rect 14606 7098 14662 7100
rect 14686 7098 14742 7100
rect 14766 7098 14822 7100
rect 14526 7046 14572 7098
rect 14572 7046 14582 7098
rect 14606 7046 14636 7098
rect 14636 7046 14648 7098
rect 14648 7046 14662 7098
rect 14686 7046 14700 7098
rect 14700 7046 14712 7098
rect 14712 7046 14742 7098
rect 14766 7046 14776 7098
rect 14776 7046 14822 7098
rect 14526 7044 14582 7046
rect 14606 7044 14662 7046
rect 14686 7044 14742 7046
rect 14766 7044 14822 7046
rect 9758 6554 9814 6556
rect 9838 6554 9894 6556
rect 9918 6554 9974 6556
rect 9998 6554 10054 6556
rect 9758 6502 9804 6554
rect 9804 6502 9814 6554
rect 9838 6502 9868 6554
rect 9868 6502 9880 6554
rect 9880 6502 9894 6554
rect 9918 6502 9932 6554
rect 9932 6502 9944 6554
rect 9944 6502 9974 6554
rect 9998 6502 10008 6554
rect 10008 6502 10054 6554
rect 9758 6500 9814 6502
rect 9838 6500 9894 6502
rect 9918 6500 9974 6502
rect 9998 6500 10054 6502
rect 15186 6554 15242 6556
rect 15266 6554 15322 6556
rect 15346 6554 15402 6556
rect 15426 6554 15482 6556
rect 15186 6502 15232 6554
rect 15232 6502 15242 6554
rect 15266 6502 15296 6554
rect 15296 6502 15308 6554
rect 15308 6502 15322 6554
rect 15346 6502 15360 6554
rect 15360 6502 15372 6554
rect 15372 6502 15402 6554
rect 15426 6502 15436 6554
rect 15436 6502 15482 6554
rect 15186 6500 15242 6502
rect 15266 6500 15322 6502
rect 15346 6500 15402 6502
rect 15426 6500 15482 6502
rect 9098 6010 9154 6012
rect 9178 6010 9234 6012
rect 9258 6010 9314 6012
rect 9338 6010 9394 6012
rect 9098 5958 9144 6010
rect 9144 5958 9154 6010
rect 9178 5958 9208 6010
rect 9208 5958 9220 6010
rect 9220 5958 9234 6010
rect 9258 5958 9272 6010
rect 9272 5958 9284 6010
rect 9284 5958 9314 6010
rect 9338 5958 9348 6010
rect 9348 5958 9394 6010
rect 9098 5956 9154 5958
rect 9178 5956 9234 5958
rect 9258 5956 9314 5958
rect 9338 5956 9394 5958
rect 14526 6010 14582 6012
rect 14606 6010 14662 6012
rect 14686 6010 14742 6012
rect 14766 6010 14822 6012
rect 14526 5958 14572 6010
rect 14572 5958 14582 6010
rect 14606 5958 14636 6010
rect 14636 5958 14648 6010
rect 14648 5958 14662 6010
rect 14686 5958 14700 6010
rect 14700 5958 14712 6010
rect 14712 5958 14742 6010
rect 14766 5958 14776 6010
rect 14776 5958 14822 6010
rect 14526 5956 14582 5958
rect 14606 5956 14662 5958
rect 14686 5956 14742 5958
rect 14766 5956 14822 5958
rect 9758 5466 9814 5468
rect 9838 5466 9894 5468
rect 9918 5466 9974 5468
rect 9998 5466 10054 5468
rect 9758 5414 9804 5466
rect 9804 5414 9814 5466
rect 9838 5414 9868 5466
rect 9868 5414 9880 5466
rect 9880 5414 9894 5466
rect 9918 5414 9932 5466
rect 9932 5414 9944 5466
rect 9944 5414 9974 5466
rect 9998 5414 10008 5466
rect 10008 5414 10054 5466
rect 9758 5412 9814 5414
rect 9838 5412 9894 5414
rect 9918 5412 9974 5414
rect 9998 5412 10054 5414
rect 15186 5466 15242 5468
rect 15266 5466 15322 5468
rect 15346 5466 15402 5468
rect 15426 5466 15482 5468
rect 15186 5414 15232 5466
rect 15232 5414 15242 5466
rect 15266 5414 15296 5466
rect 15296 5414 15308 5466
rect 15308 5414 15322 5466
rect 15346 5414 15360 5466
rect 15360 5414 15372 5466
rect 15372 5414 15402 5466
rect 15426 5414 15436 5466
rect 15436 5414 15482 5466
rect 15186 5412 15242 5414
rect 15266 5412 15322 5414
rect 15346 5412 15402 5414
rect 15426 5412 15482 5414
rect 9098 4922 9154 4924
rect 9178 4922 9234 4924
rect 9258 4922 9314 4924
rect 9338 4922 9394 4924
rect 9098 4870 9144 4922
rect 9144 4870 9154 4922
rect 9178 4870 9208 4922
rect 9208 4870 9220 4922
rect 9220 4870 9234 4922
rect 9258 4870 9272 4922
rect 9272 4870 9284 4922
rect 9284 4870 9314 4922
rect 9338 4870 9348 4922
rect 9348 4870 9394 4922
rect 9098 4868 9154 4870
rect 9178 4868 9234 4870
rect 9258 4868 9314 4870
rect 9338 4868 9394 4870
rect 14526 4922 14582 4924
rect 14606 4922 14662 4924
rect 14686 4922 14742 4924
rect 14766 4922 14822 4924
rect 14526 4870 14572 4922
rect 14572 4870 14582 4922
rect 14606 4870 14636 4922
rect 14636 4870 14648 4922
rect 14648 4870 14662 4922
rect 14686 4870 14700 4922
rect 14700 4870 14712 4922
rect 14712 4870 14742 4922
rect 14766 4870 14776 4922
rect 14776 4870 14822 4922
rect 14526 4868 14582 4870
rect 14606 4868 14662 4870
rect 14686 4868 14742 4870
rect 14766 4868 14822 4870
rect 9758 4378 9814 4380
rect 9838 4378 9894 4380
rect 9918 4378 9974 4380
rect 9998 4378 10054 4380
rect 9758 4326 9804 4378
rect 9804 4326 9814 4378
rect 9838 4326 9868 4378
rect 9868 4326 9880 4378
rect 9880 4326 9894 4378
rect 9918 4326 9932 4378
rect 9932 4326 9944 4378
rect 9944 4326 9974 4378
rect 9998 4326 10008 4378
rect 10008 4326 10054 4378
rect 9758 4324 9814 4326
rect 9838 4324 9894 4326
rect 9918 4324 9974 4326
rect 9998 4324 10054 4326
rect 15186 4378 15242 4380
rect 15266 4378 15322 4380
rect 15346 4378 15402 4380
rect 15426 4378 15482 4380
rect 15186 4326 15232 4378
rect 15232 4326 15242 4378
rect 15266 4326 15296 4378
rect 15296 4326 15308 4378
rect 15308 4326 15322 4378
rect 15346 4326 15360 4378
rect 15360 4326 15372 4378
rect 15372 4326 15402 4378
rect 15426 4326 15436 4378
rect 15436 4326 15482 4378
rect 15186 4324 15242 4326
rect 15266 4324 15322 4326
rect 15346 4324 15402 4326
rect 15426 4324 15482 4326
rect 3670 3834 3726 3836
rect 3750 3834 3806 3836
rect 3830 3834 3886 3836
rect 3910 3834 3966 3836
rect 3670 3782 3716 3834
rect 3716 3782 3726 3834
rect 3750 3782 3780 3834
rect 3780 3782 3792 3834
rect 3792 3782 3806 3834
rect 3830 3782 3844 3834
rect 3844 3782 3856 3834
rect 3856 3782 3886 3834
rect 3910 3782 3920 3834
rect 3920 3782 3966 3834
rect 3670 3780 3726 3782
rect 3750 3780 3806 3782
rect 3830 3780 3886 3782
rect 3910 3780 3966 3782
rect 4330 3290 4386 3292
rect 4410 3290 4466 3292
rect 4490 3290 4546 3292
rect 4570 3290 4626 3292
rect 4330 3238 4376 3290
rect 4376 3238 4386 3290
rect 4410 3238 4440 3290
rect 4440 3238 4452 3290
rect 4452 3238 4466 3290
rect 4490 3238 4504 3290
rect 4504 3238 4516 3290
rect 4516 3238 4546 3290
rect 4570 3238 4580 3290
rect 4580 3238 4626 3290
rect 4330 3236 4386 3238
rect 4410 3236 4466 3238
rect 4490 3236 4546 3238
rect 4570 3236 4626 3238
rect 3670 2746 3726 2748
rect 3750 2746 3806 2748
rect 3830 2746 3886 2748
rect 3910 2746 3966 2748
rect 3670 2694 3716 2746
rect 3716 2694 3726 2746
rect 3750 2694 3780 2746
rect 3780 2694 3792 2746
rect 3792 2694 3806 2746
rect 3830 2694 3844 2746
rect 3844 2694 3856 2746
rect 3856 2694 3886 2746
rect 3910 2694 3920 2746
rect 3920 2694 3966 2746
rect 3670 2692 3726 2694
rect 3750 2692 3806 2694
rect 3830 2692 3886 2694
rect 3910 2692 3966 2694
rect 9098 3834 9154 3836
rect 9178 3834 9234 3836
rect 9258 3834 9314 3836
rect 9338 3834 9394 3836
rect 9098 3782 9144 3834
rect 9144 3782 9154 3834
rect 9178 3782 9208 3834
rect 9208 3782 9220 3834
rect 9220 3782 9234 3834
rect 9258 3782 9272 3834
rect 9272 3782 9284 3834
rect 9284 3782 9314 3834
rect 9338 3782 9348 3834
rect 9348 3782 9394 3834
rect 9098 3780 9154 3782
rect 9178 3780 9234 3782
rect 9258 3780 9314 3782
rect 9338 3780 9394 3782
rect 14526 3834 14582 3836
rect 14606 3834 14662 3836
rect 14686 3834 14742 3836
rect 14766 3834 14822 3836
rect 14526 3782 14572 3834
rect 14572 3782 14582 3834
rect 14606 3782 14636 3834
rect 14636 3782 14648 3834
rect 14648 3782 14662 3834
rect 14686 3782 14700 3834
rect 14700 3782 14712 3834
rect 14712 3782 14742 3834
rect 14766 3782 14776 3834
rect 14776 3782 14822 3834
rect 14526 3780 14582 3782
rect 14606 3780 14662 3782
rect 14686 3780 14742 3782
rect 14766 3780 14822 3782
rect 9758 3290 9814 3292
rect 9838 3290 9894 3292
rect 9918 3290 9974 3292
rect 9998 3290 10054 3292
rect 9758 3238 9804 3290
rect 9804 3238 9814 3290
rect 9838 3238 9868 3290
rect 9868 3238 9880 3290
rect 9880 3238 9894 3290
rect 9918 3238 9932 3290
rect 9932 3238 9944 3290
rect 9944 3238 9974 3290
rect 9998 3238 10008 3290
rect 10008 3238 10054 3290
rect 9758 3236 9814 3238
rect 9838 3236 9894 3238
rect 9918 3236 9974 3238
rect 9998 3236 10054 3238
rect 15186 3290 15242 3292
rect 15266 3290 15322 3292
rect 15346 3290 15402 3292
rect 15426 3290 15482 3292
rect 15186 3238 15232 3290
rect 15232 3238 15242 3290
rect 15266 3238 15296 3290
rect 15296 3238 15308 3290
rect 15308 3238 15322 3290
rect 15346 3238 15360 3290
rect 15360 3238 15372 3290
rect 15372 3238 15402 3290
rect 15426 3238 15436 3290
rect 15436 3238 15482 3290
rect 15186 3236 15242 3238
rect 15266 3236 15322 3238
rect 15346 3236 15402 3238
rect 15426 3236 15482 3238
rect 9098 2746 9154 2748
rect 9178 2746 9234 2748
rect 9258 2746 9314 2748
rect 9338 2746 9394 2748
rect 9098 2694 9144 2746
rect 9144 2694 9154 2746
rect 9178 2694 9208 2746
rect 9208 2694 9220 2746
rect 9220 2694 9234 2746
rect 9258 2694 9272 2746
rect 9272 2694 9284 2746
rect 9284 2694 9314 2746
rect 9338 2694 9348 2746
rect 9348 2694 9394 2746
rect 9098 2692 9154 2694
rect 9178 2692 9234 2694
rect 9258 2692 9314 2694
rect 9338 2692 9394 2694
rect 14526 2746 14582 2748
rect 14606 2746 14662 2748
rect 14686 2746 14742 2748
rect 14766 2746 14822 2748
rect 14526 2694 14572 2746
rect 14572 2694 14582 2746
rect 14606 2694 14636 2746
rect 14636 2694 14648 2746
rect 14648 2694 14662 2746
rect 14686 2694 14700 2746
rect 14700 2694 14712 2746
rect 14712 2694 14742 2746
rect 14766 2694 14776 2746
rect 14776 2694 14822 2746
rect 14526 2692 14582 2694
rect 14606 2692 14662 2694
rect 14686 2692 14742 2694
rect 14766 2692 14822 2694
rect 20614 17434 20670 17436
rect 20694 17434 20750 17436
rect 20774 17434 20830 17436
rect 20854 17434 20910 17436
rect 20614 17382 20660 17434
rect 20660 17382 20670 17434
rect 20694 17382 20724 17434
rect 20724 17382 20736 17434
rect 20736 17382 20750 17434
rect 20774 17382 20788 17434
rect 20788 17382 20800 17434
rect 20800 17382 20830 17434
rect 20854 17382 20864 17434
rect 20864 17382 20910 17434
rect 20614 17380 20670 17382
rect 20694 17380 20750 17382
rect 20774 17380 20830 17382
rect 20854 17380 20910 17382
rect 19954 16890 20010 16892
rect 20034 16890 20090 16892
rect 20114 16890 20170 16892
rect 20194 16890 20250 16892
rect 19954 16838 20000 16890
rect 20000 16838 20010 16890
rect 20034 16838 20064 16890
rect 20064 16838 20076 16890
rect 20076 16838 20090 16890
rect 20114 16838 20128 16890
rect 20128 16838 20140 16890
rect 20140 16838 20170 16890
rect 20194 16838 20204 16890
rect 20204 16838 20250 16890
rect 19954 16836 20010 16838
rect 20034 16836 20090 16838
rect 20114 16836 20170 16838
rect 20194 16836 20250 16838
rect 20614 16346 20670 16348
rect 20694 16346 20750 16348
rect 20774 16346 20830 16348
rect 20854 16346 20910 16348
rect 20614 16294 20660 16346
rect 20660 16294 20670 16346
rect 20694 16294 20724 16346
rect 20724 16294 20736 16346
rect 20736 16294 20750 16346
rect 20774 16294 20788 16346
rect 20788 16294 20800 16346
rect 20800 16294 20830 16346
rect 20854 16294 20864 16346
rect 20864 16294 20910 16346
rect 20614 16292 20670 16294
rect 20694 16292 20750 16294
rect 20774 16292 20830 16294
rect 20854 16292 20910 16294
rect 19954 15802 20010 15804
rect 20034 15802 20090 15804
rect 20114 15802 20170 15804
rect 20194 15802 20250 15804
rect 19954 15750 20000 15802
rect 20000 15750 20010 15802
rect 20034 15750 20064 15802
rect 20064 15750 20076 15802
rect 20076 15750 20090 15802
rect 20114 15750 20128 15802
rect 20128 15750 20140 15802
rect 20140 15750 20170 15802
rect 20194 15750 20204 15802
rect 20204 15750 20250 15802
rect 19954 15748 20010 15750
rect 20034 15748 20090 15750
rect 20114 15748 20170 15750
rect 20194 15748 20250 15750
rect 20614 15258 20670 15260
rect 20694 15258 20750 15260
rect 20774 15258 20830 15260
rect 20854 15258 20910 15260
rect 20614 15206 20660 15258
rect 20660 15206 20670 15258
rect 20694 15206 20724 15258
rect 20724 15206 20736 15258
rect 20736 15206 20750 15258
rect 20774 15206 20788 15258
rect 20788 15206 20800 15258
rect 20800 15206 20830 15258
rect 20854 15206 20864 15258
rect 20864 15206 20910 15258
rect 20614 15204 20670 15206
rect 20694 15204 20750 15206
rect 20774 15204 20830 15206
rect 20854 15204 20910 15206
rect 19954 14714 20010 14716
rect 20034 14714 20090 14716
rect 20114 14714 20170 14716
rect 20194 14714 20250 14716
rect 19954 14662 20000 14714
rect 20000 14662 20010 14714
rect 20034 14662 20064 14714
rect 20064 14662 20076 14714
rect 20076 14662 20090 14714
rect 20114 14662 20128 14714
rect 20128 14662 20140 14714
rect 20140 14662 20170 14714
rect 20194 14662 20204 14714
rect 20204 14662 20250 14714
rect 19954 14660 20010 14662
rect 20034 14660 20090 14662
rect 20114 14660 20170 14662
rect 20194 14660 20250 14662
rect 20614 14170 20670 14172
rect 20694 14170 20750 14172
rect 20774 14170 20830 14172
rect 20854 14170 20910 14172
rect 20614 14118 20660 14170
rect 20660 14118 20670 14170
rect 20694 14118 20724 14170
rect 20724 14118 20736 14170
rect 20736 14118 20750 14170
rect 20774 14118 20788 14170
rect 20788 14118 20800 14170
rect 20800 14118 20830 14170
rect 20854 14118 20864 14170
rect 20864 14118 20910 14170
rect 20614 14116 20670 14118
rect 20694 14116 20750 14118
rect 20774 14116 20830 14118
rect 20854 14116 20910 14118
rect 19954 13626 20010 13628
rect 20034 13626 20090 13628
rect 20114 13626 20170 13628
rect 20194 13626 20250 13628
rect 19954 13574 20000 13626
rect 20000 13574 20010 13626
rect 20034 13574 20064 13626
rect 20064 13574 20076 13626
rect 20076 13574 20090 13626
rect 20114 13574 20128 13626
rect 20128 13574 20140 13626
rect 20140 13574 20170 13626
rect 20194 13574 20204 13626
rect 20204 13574 20250 13626
rect 19954 13572 20010 13574
rect 20034 13572 20090 13574
rect 20114 13572 20170 13574
rect 20194 13572 20250 13574
rect 20614 13082 20670 13084
rect 20694 13082 20750 13084
rect 20774 13082 20830 13084
rect 20854 13082 20910 13084
rect 20614 13030 20660 13082
rect 20660 13030 20670 13082
rect 20694 13030 20724 13082
rect 20724 13030 20736 13082
rect 20736 13030 20750 13082
rect 20774 13030 20788 13082
rect 20788 13030 20800 13082
rect 20800 13030 20830 13082
rect 20854 13030 20864 13082
rect 20864 13030 20910 13082
rect 20614 13028 20670 13030
rect 20694 13028 20750 13030
rect 20774 13028 20830 13030
rect 20854 13028 20910 13030
rect 19954 12538 20010 12540
rect 20034 12538 20090 12540
rect 20114 12538 20170 12540
rect 20194 12538 20250 12540
rect 19954 12486 20000 12538
rect 20000 12486 20010 12538
rect 20034 12486 20064 12538
rect 20064 12486 20076 12538
rect 20076 12486 20090 12538
rect 20114 12486 20128 12538
rect 20128 12486 20140 12538
rect 20140 12486 20170 12538
rect 20194 12486 20204 12538
rect 20204 12486 20250 12538
rect 19954 12484 20010 12486
rect 20034 12484 20090 12486
rect 20114 12484 20170 12486
rect 20194 12484 20250 12486
rect 20614 11994 20670 11996
rect 20694 11994 20750 11996
rect 20774 11994 20830 11996
rect 20854 11994 20910 11996
rect 20614 11942 20660 11994
rect 20660 11942 20670 11994
rect 20694 11942 20724 11994
rect 20724 11942 20736 11994
rect 20736 11942 20750 11994
rect 20774 11942 20788 11994
rect 20788 11942 20800 11994
rect 20800 11942 20830 11994
rect 20854 11942 20864 11994
rect 20864 11942 20910 11994
rect 20614 11940 20670 11942
rect 20694 11940 20750 11942
rect 20774 11940 20830 11942
rect 20854 11940 20910 11942
rect 19954 11450 20010 11452
rect 20034 11450 20090 11452
rect 20114 11450 20170 11452
rect 20194 11450 20250 11452
rect 19954 11398 20000 11450
rect 20000 11398 20010 11450
rect 20034 11398 20064 11450
rect 20064 11398 20076 11450
rect 20076 11398 20090 11450
rect 20114 11398 20128 11450
rect 20128 11398 20140 11450
rect 20140 11398 20170 11450
rect 20194 11398 20204 11450
rect 20204 11398 20250 11450
rect 19954 11396 20010 11398
rect 20034 11396 20090 11398
rect 20114 11396 20170 11398
rect 20194 11396 20250 11398
rect 20614 10906 20670 10908
rect 20694 10906 20750 10908
rect 20774 10906 20830 10908
rect 20854 10906 20910 10908
rect 20614 10854 20660 10906
rect 20660 10854 20670 10906
rect 20694 10854 20724 10906
rect 20724 10854 20736 10906
rect 20736 10854 20750 10906
rect 20774 10854 20788 10906
rect 20788 10854 20800 10906
rect 20800 10854 20830 10906
rect 20854 10854 20864 10906
rect 20864 10854 20910 10906
rect 20614 10852 20670 10854
rect 20694 10852 20750 10854
rect 20774 10852 20830 10854
rect 20854 10852 20910 10854
rect 19954 10362 20010 10364
rect 20034 10362 20090 10364
rect 20114 10362 20170 10364
rect 20194 10362 20250 10364
rect 19954 10310 20000 10362
rect 20000 10310 20010 10362
rect 20034 10310 20064 10362
rect 20064 10310 20076 10362
rect 20076 10310 20090 10362
rect 20114 10310 20128 10362
rect 20128 10310 20140 10362
rect 20140 10310 20170 10362
rect 20194 10310 20204 10362
rect 20204 10310 20250 10362
rect 19954 10308 20010 10310
rect 20034 10308 20090 10310
rect 20114 10308 20170 10310
rect 20194 10308 20250 10310
rect 22374 10240 22430 10296
rect 20614 9818 20670 9820
rect 20694 9818 20750 9820
rect 20774 9818 20830 9820
rect 20854 9818 20910 9820
rect 20614 9766 20660 9818
rect 20660 9766 20670 9818
rect 20694 9766 20724 9818
rect 20724 9766 20736 9818
rect 20736 9766 20750 9818
rect 20774 9766 20788 9818
rect 20788 9766 20800 9818
rect 20800 9766 20830 9818
rect 20854 9766 20864 9818
rect 20864 9766 20910 9818
rect 20614 9764 20670 9766
rect 20694 9764 20750 9766
rect 20774 9764 20830 9766
rect 20854 9764 20910 9766
rect 19954 9274 20010 9276
rect 20034 9274 20090 9276
rect 20114 9274 20170 9276
rect 20194 9274 20250 9276
rect 19954 9222 20000 9274
rect 20000 9222 20010 9274
rect 20034 9222 20064 9274
rect 20064 9222 20076 9274
rect 20076 9222 20090 9274
rect 20114 9222 20128 9274
rect 20128 9222 20140 9274
rect 20140 9222 20170 9274
rect 20194 9222 20204 9274
rect 20204 9222 20250 9274
rect 19954 9220 20010 9222
rect 20034 9220 20090 9222
rect 20114 9220 20170 9222
rect 20194 9220 20250 9222
rect 20614 8730 20670 8732
rect 20694 8730 20750 8732
rect 20774 8730 20830 8732
rect 20854 8730 20910 8732
rect 20614 8678 20660 8730
rect 20660 8678 20670 8730
rect 20694 8678 20724 8730
rect 20724 8678 20736 8730
rect 20736 8678 20750 8730
rect 20774 8678 20788 8730
rect 20788 8678 20800 8730
rect 20800 8678 20830 8730
rect 20854 8678 20864 8730
rect 20864 8678 20910 8730
rect 20614 8676 20670 8678
rect 20694 8676 20750 8678
rect 20774 8676 20830 8678
rect 20854 8676 20910 8678
rect 19954 8186 20010 8188
rect 20034 8186 20090 8188
rect 20114 8186 20170 8188
rect 20194 8186 20250 8188
rect 19954 8134 20000 8186
rect 20000 8134 20010 8186
rect 20034 8134 20064 8186
rect 20064 8134 20076 8186
rect 20076 8134 20090 8186
rect 20114 8134 20128 8186
rect 20128 8134 20140 8186
rect 20140 8134 20170 8186
rect 20194 8134 20204 8186
rect 20204 8134 20250 8186
rect 19954 8132 20010 8134
rect 20034 8132 20090 8134
rect 20114 8132 20170 8134
rect 20194 8132 20250 8134
rect 20614 7642 20670 7644
rect 20694 7642 20750 7644
rect 20774 7642 20830 7644
rect 20854 7642 20910 7644
rect 20614 7590 20660 7642
rect 20660 7590 20670 7642
rect 20694 7590 20724 7642
rect 20724 7590 20736 7642
rect 20736 7590 20750 7642
rect 20774 7590 20788 7642
rect 20788 7590 20800 7642
rect 20800 7590 20830 7642
rect 20854 7590 20864 7642
rect 20864 7590 20910 7642
rect 20614 7588 20670 7590
rect 20694 7588 20750 7590
rect 20774 7588 20830 7590
rect 20854 7588 20910 7590
rect 19954 7098 20010 7100
rect 20034 7098 20090 7100
rect 20114 7098 20170 7100
rect 20194 7098 20250 7100
rect 19954 7046 20000 7098
rect 20000 7046 20010 7098
rect 20034 7046 20064 7098
rect 20064 7046 20076 7098
rect 20076 7046 20090 7098
rect 20114 7046 20128 7098
rect 20128 7046 20140 7098
rect 20140 7046 20170 7098
rect 20194 7046 20204 7098
rect 20204 7046 20250 7098
rect 19954 7044 20010 7046
rect 20034 7044 20090 7046
rect 20114 7044 20170 7046
rect 20194 7044 20250 7046
rect 20614 6554 20670 6556
rect 20694 6554 20750 6556
rect 20774 6554 20830 6556
rect 20854 6554 20910 6556
rect 20614 6502 20660 6554
rect 20660 6502 20670 6554
rect 20694 6502 20724 6554
rect 20724 6502 20736 6554
rect 20736 6502 20750 6554
rect 20774 6502 20788 6554
rect 20788 6502 20800 6554
rect 20800 6502 20830 6554
rect 20854 6502 20864 6554
rect 20864 6502 20910 6554
rect 20614 6500 20670 6502
rect 20694 6500 20750 6502
rect 20774 6500 20830 6502
rect 20854 6500 20910 6502
rect 19954 6010 20010 6012
rect 20034 6010 20090 6012
rect 20114 6010 20170 6012
rect 20194 6010 20250 6012
rect 19954 5958 20000 6010
rect 20000 5958 20010 6010
rect 20034 5958 20064 6010
rect 20064 5958 20076 6010
rect 20076 5958 20090 6010
rect 20114 5958 20128 6010
rect 20128 5958 20140 6010
rect 20140 5958 20170 6010
rect 20194 5958 20204 6010
rect 20204 5958 20250 6010
rect 19954 5956 20010 5958
rect 20034 5956 20090 5958
rect 20114 5956 20170 5958
rect 20194 5956 20250 5958
rect 20614 5466 20670 5468
rect 20694 5466 20750 5468
rect 20774 5466 20830 5468
rect 20854 5466 20910 5468
rect 20614 5414 20660 5466
rect 20660 5414 20670 5466
rect 20694 5414 20724 5466
rect 20724 5414 20736 5466
rect 20736 5414 20750 5466
rect 20774 5414 20788 5466
rect 20788 5414 20800 5466
rect 20800 5414 20830 5466
rect 20854 5414 20864 5466
rect 20864 5414 20910 5466
rect 20614 5412 20670 5414
rect 20694 5412 20750 5414
rect 20774 5412 20830 5414
rect 20854 5412 20910 5414
rect 19954 4922 20010 4924
rect 20034 4922 20090 4924
rect 20114 4922 20170 4924
rect 20194 4922 20250 4924
rect 19954 4870 20000 4922
rect 20000 4870 20010 4922
rect 20034 4870 20064 4922
rect 20064 4870 20076 4922
rect 20076 4870 20090 4922
rect 20114 4870 20128 4922
rect 20128 4870 20140 4922
rect 20140 4870 20170 4922
rect 20194 4870 20204 4922
rect 20204 4870 20250 4922
rect 19954 4868 20010 4870
rect 20034 4868 20090 4870
rect 20114 4868 20170 4870
rect 20194 4868 20250 4870
rect 20614 4378 20670 4380
rect 20694 4378 20750 4380
rect 20774 4378 20830 4380
rect 20854 4378 20910 4380
rect 20614 4326 20660 4378
rect 20660 4326 20670 4378
rect 20694 4326 20724 4378
rect 20724 4326 20736 4378
rect 20736 4326 20750 4378
rect 20774 4326 20788 4378
rect 20788 4326 20800 4378
rect 20800 4326 20830 4378
rect 20854 4326 20864 4378
rect 20864 4326 20910 4378
rect 20614 4324 20670 4326
rect 20694 4324 20750 4326
rect 20774 4324 20830 4326
rect 20854 4324 20910 4326
rect 19954 3834 20010 3836
rect 20034 3834 20090 3836
rect 20114 3834 20170 3836
rect 20194 3834 20250 3836
rect 19954 3782 20000 3834
rect 20000 3782 20010 3834
rect 20034 3782 20064 3834
rect 20064 3782 20076 3834
rect 20076 3782 20090 3834
rect 20114 3782 20128 3834
rect 20128 3782 20140 3834
rect 20140 3782 20170 3834
rect 20194 3782 20204 3834
rect 20204 3782 20250 3834
rect 19954 3780 20010 3782
rect 20034 3780 20090 3782
rect 20114 3780 20170 3782
rect 20194 3780 20250 3782
rect 20614 3290 20670 3292
rect 20694 3290 20750 3292
rect 20774 3290 20830 3292
rect 20854 3290 20910 3292
rect 20614 3238 20660 3290
rect 20660 3238 20670 3290
rect 20694 3238 20724 3290
rect 20724 3238 20736 3290
rect 20736 3238 20750 3290
rect 20774 3238 20788 3290
rect 20788 3238 20800 3290
rect 20800 3238 20830 3290
rect 20854 3238 20864 3290
rect 20864 3238 20910 3290
rect 20614 3236 20670 3238
rect 20694 3236 20750 3238
rect 20774 3236 20830 3238
rect 20854 3236 20910 3238
rect 19954 2746 20010 2748
rect 20034 2746 20090 2748
rect 20114 2746 20170 2748
rect 20194 2746 20250 2748
rect 19954 2694 20000 2746
rect 20000 2694 20010 2746
rect 20034 2694 20064 2746
rect 20064 2694 20076 2746
rect 20076 2694 20090 2746
rect 20114 2694 20128 2746
rect 20128 2694 20140 2746
rect 20140 2694 20170 2746
rect 20194 2694 20204 2746
rect 20204 2694 20250 2746
rect 19954 2692 20010 2694
rect 20034 2692 20090 2694
rect 20114 2692 20170 2694
rect 20194 2692 20250 2694
rect 4330 2202 4386 2204
rect 4410 2202 4466 2204
rect 4490 2202 4546 2204
rect 4570 2202 4626 2204
rect 4330 2150 4376 2202
rect 4376 2150 4386 2202
rect 4410 2150 4440 2202
rect 4440 2150 4452 2202
rect 4452 2150 4466 2202
rect 4490 2150 4504 2202
rect 4504 2150 4516 2202
rect 4516 2150 4546 2202
rect 4570 2150 4580 2202
rect 4580 2150 4626 2202
rect 4330 2148 4386 2150
rect 4410 2148 4466 2150
rect 4490 2148 4546 2150
rect 4570 2148 4626 2150
rect 9758 2202 9814 2204
rect 9838 2202 9894 2204
rect 9918 2202 9974 2204
rect 9998 2202 10054 2204
rect 9758 2150 9804 2202
rect 9804 2150 9814 2202
rect 9838 2150 9868 2202
rect 9868 2150 9880 2202
rect 9880 2150 9894 2202
rect 9918 2150 9932 2202
rect 9932 2150 9944 2202
rect 9944 2150 9974 2202
rect 9998 2150 10008 2202
rect 10008 2150 10054 2202
rect 9758 2148 9814 2150
rect 9838 2148 9894 2150
rect 9918 2148 9974 2150
rect 9998 2148 10054 2150
rect 15186 2202 15242 2204
rect 15266 2202 15322 2204
rect 15346 2202 15402 2204
rect 15426 2202 15482 2204
rect 15186 2150 15232 2202
rect 15232 2150 15242 2202
rect 15266 2150 15296 2202
rect 15296 2150 15308 2202
rect 15308 2150 15322 2202
rect 15346 2150 15360 2202
rect 15360 2150 15372 2202
rect 15372 2150 15402 2202
rect 15426 2150 15436 2202
rect 15436 2150 15482 2202
rect 15186 2148 15242 2150
rect 15266 2148 15322 2150
rect 15346 2148 15402 2150
rect 15426 2148 15482 2150
rect 20614 2202 20670 2204
rect 20694 2202 20750 2204
rect 20774 2202 20830 2204
rect 20854 2202 20910 2204
rect 20614 2150 20660 2202
rect 20660 2150 20670 2202
rect 20694 2150 20724 2202
rect 20724 2150 20736 2202
rect 20736 2150 20750 2202
rect 20774 2150 20788 2202
rect 20788 2150 20800 2202
rect 20800 2150 20830 2202
rect 20854 2150 20864 2202
rect 20864 2150 20910 2202
rect 20614 2148 20670 2150
rect 20694 2148 20750 2150
rect 20774 2148 20830 2150
rect 20854 2148 20910 2150
rect 22834 1400 22890 1456
<< metal3 >>
rect 4320 21792 4636 21793
rect 4320 21728 4326 21792
rect 4390 21728 4406 21792
rect 4470 21728 4486 21792
rect 4550 21728 4566 21792
rect 4630 21728 4636 21792
rect 4320 21727 4636 21728
rect 9748 21792 10064 21793
rect 9748 21728 9754 21792
rect 9818 21728 9834 21792
rect 9898 21728 9914 21792
rect 9978 21728 9994 21792
rect 10058 21728 10064 21792
rect 9748 21727 10064 21728
rect 15176 21792 15492 21793
rect 15176 21728 15182 21792
rect 15246 21728 15262 21792
rect 15326 21728 15342 21792
rect 15406 21728 15422 21792
rect 15486 21728 15492 21792
rect 15176 21727 15492 21728
rect 20604 21792 20920 21793
rect 20604 21728 20610 21792
rect 20674 21728 20690 21792
rect 20754 21728 20770 21792
rect 20834 21728 20850 21792
rect 20914 21728 20920 21792
rect 20604 21727 20920 21728
rect 3660 21248 3976 21249
rect 3660 21184 3666 21248
rect 3730 21184 3746 21248
rect 3810 21184 3826 21248
rect 3890 21184 3906 21248
rect 3970 21184 3976 21248
rect 3660 21183 3976 21184
rect 9088 21248 9404 21249
rect 9088 21184 9094 21248
rect 9158 21184 9174 21248
rect 9238 21184 9254 21248
rect 9318 21184 9334 21248
rect 9398 21184 9404 21248
rect 9088 21183 9404 21184
rect 14516 21248 14832 21249
rect 14516 21184 14522 21248
rect 14586 21184 14602 21248
rect 14666 21184 14682 21248
rect 14746 21184 14762 21248
rect 14826 21184 14832 21248
rect 14516 21183 14832 21184
rect 19944 21248 20260 21249
rect 19944 21184 19950 21248
rect 20014 21184 20030 21248
rect 20094 21184 20110 21248
rect 20174 21184 20190 21248
rect 20254 21184 20260 21248
rect 19944 21183 20260 21184
rect 4320 20704 4636 20705
rect 4320 20640 4326 20704
rect 4390 20640 4406 20704
rect 4470 20640 4486 20704
rect 4550 20640 4566 20704
rect 4630 20640 4636 20704
rect 4320 20639 4636 20640
rect 9748 20704 10064 20705
rect 9748 20640 9754 20704
rect 9818 20640 9834 20704
rect 9898 20640 9914 20704
rect 9978 20640 9994 20704
rect 10058 20640 10064 20704
rect 9748 20639 10064 20640
rect 15176 20704 15492 20705
rect 15176 20640 15182 20704
rect 15246 20640 15262 20704
rect 15326 20640 15342 20704
rect 15406 20640 15422 20704
rect 15486 20640 15492 20704
rect 15176 20639 15492 20640
rect 20604 20704 20920 20705
rect 20604 20640 20610 20704
rect 20674 20640 20690 20704
rect 20754 20640 20770 20704
rect 20834 20640 20850 20704
rect 20914 20640 20920 20704
rect 20604 20639 20920 20640
rect 3660 20160 3976 20161
rect 3660 20096 3666 20160
rect 3730 20096 3746 20160
rect 3810 20096 3826 20160
rect 3890 20096 3906 20160
rect 3970 20096 3976 20160
rect 3660 20095 3976 20096
rect 9088 20160 9404 20161
rect 9088 20096 9094 20160
rect 9158 20096 9174 20160
rect 9238 20096 9254 20160
rect 9318 20096 9334 20160
rect 9398 20096 9404 20160
rect 9088 20095 9404 20096
rect 14516 20160 14832 20161
rect 14516 20096 14522 20160
rect 14586 20096 14602 20160
rect 14666 20096 14682 20160
rect 14746 20096 14762 20160
rect 14826 20096 14832 20160
rect 14516 20095 14832 20096
rect 19944 20160 20260 20161
rect 19944 20096 19950 20160
rect 20014 20096 20030 20160
rect 20094 20096 20110 20160
rect 20174 20096 20190 20160
rect 20254 20096 20260 20160
rect 19944 20095 20260 20096
rect 22829 19818 22895 19821
rect 23200 19818 24000 19848
rect 22829 19816 24000 19818
rect 22829 19760 22834 19816
rect 22890 19760 24000 19816
rect 22829 19758 24000 19760
rect 22829 19755 22895 19758
rect 23200 19728 24000 19758
rect 4320 19616 4636 19617
rect 4320 19552 4326 19616
rect 4390 19552 4406 19616
rect 4470 19552 4486 19616
rect 4550 19552 4566 19616
rect 4630 19552 4636 19616
rect 4320 19551 4636 19552
rect 9748 19616 10064 19617
rect 9748 19552 9754 19616
rect 9818 19552 9834 19616
rect 9898 19552 9914 19616
rect 9978 19552 9994 19616
rect 10058 19552 10064 19616
rect 9748 19551 10064 19552
rect 15176 19616 15492 19617
rect 15176 19552 15182 19616
rect 15246 19552 15262 19616
rect 15326 19552 15342 19616
rect 15406 19552 15422 19616
rect 15486 19552 15492 19616
rect 15176 19551 15492 19552
rect 20604 19616 20920 19617
rect 20604 19552 20610 19616
rect 20674 19552 20690 19616
rect 20754 19552 20770 19616
rect 20834 19552 20850 19616
rect 20914 19552 20920 19616
rect 20604 19551 20920 19552
rect 3660 19072 3976 19073
rect 3660 19008 3666 19072
rect 3730 19008 3746 19072
rect 3810 19008 3826 19072
rect 3890 19008 3906 19072
rect 3970 19008 3976 19072
rect 3660 19007 3976 19008
rect 9088 19072 9404 19073
rect 9088 19008 9094 19072
rect 9158 19008 9174 19072
rect 9238 19008 9254 19072
rect 9318 19008 9334 19072
rect 9398 19008 9404 19072
rect 9088 19007 9404 19008
rect 14516 19072 14832 19073
rect 14516 19008 14522 19072
rect 14586 19008 14602 19072
rect 14666 19008 14682 19072
rect 14746 19008 14762 19072
rect 14826 19008 14832 19072
rect 14516 19007 14832 19008
rect 19944 19072 20260 19073
rect 19944 19008 19950 19072
rect 20014 19008 20030 19072
rect 20094 19008 20110 19072
rect 20174 19008 20190 19072
rect 20254 19008 20260 19072
rect 19944 19007 20260 19008
rect 4320 18528 4636 18529
rect 4320 18464 4326 18528
rect 4390 18464 4406 18528
rect 4470 18464 4486 18528
rect 4550 18464 4566 18528
rect 4630 18464 4636 18528
rect 4320 18463 4636 18464
rect 9748 18528 10064 18529
rect 9748 18464 9754 18528
rect 9818 18464 9834 18528
rect 9898 18464 9914 18528
rect 9978 18464 9994 18528
rect 10058 18464 10064 18528
rect 9748 18463 10064 18464
rect 15176 18528 15492 18529
rect 15176 18464 15182 18528
rect 15246 18464 15262 18528
rect 15326 18464 15342 18528
rect 15406 18464 15422 18528
rect 15486 18464 15492 18528
rect 15176 18463 15492 18464
rect 20604 18528 20920 18529
rect 20604 18464 20610 18528
rect 20674 18464 20690 18528
rect 20754 18464 20770 18528
rect 20834 18464 20850 18528
rect 20914 18464 20920 18528
rect 20604 18463 20920 18464
rect 3660 17984 3976 17985
rect 3660 17920 3666 17984
rect 3730 17920 3746 17984
rect 3810 17920 3826 17984
rect 3890 17920 3906 17984
rect 3970 17920 3976 17984
rect 3660 17919 3976 17920
rect 9088 17984 9404 17985
rect 9088 17920 9094 17984
rect 9158 17920 9174 17984
rect 9238 17920 9254 17984
rect 9318 17920 9334 17984
rect 9398 17920 9404 17984
rect 9088 17919 9404 17920
rect 14516 17984 14832 17985
rect 14516 17920 14522 17984
rect 14586 17920 14602 17984
rect 14666 17920 14682 17984
rect 14746 17920 14762 17984
rect 14826 17920 14832 17984
rect 14516 17919 14832 17920
rect 19944 17984 20260 17985
rect 19944 17920 19950 17984
rect 20014 17920 20030 17984
rect 20094 17920 20110 17984
rect 20174 17920 20190 17984
rect 20254 17920 20260 17984
rect 19944 17919 20260 17920
rect 1485 17914 1551 17917
rect 798 17912 1551 17914
rect 798 17856 1490 17912
rect 1546 17856 1551 17912
rect 798 17854 1551 17856
rect 798 17808 858 17854
rect 1485 17851 1551 17854
rect 0 17718 858 17808
rect 0 17688 800 17718
rect 4320 17440 4636 17441
rect 4320 17376 4326 17440
rect 4390 17376 4406 17440
rect 4470 17376 4486 17440
rect 4550 17376 4566 17440
rect 4630 17376 4636 17440
rect 4320 17375 4636 17376
rect 9748 17440 10064 17441
rect 9748 17376 9754 17440
rect 9818 17376 9834 17440
rect 9898 17376 9914 17440
rect 9978 17376 9994 17440
rect 10058 17376 10064 17440
rect 9748 17375 10064 17376
rect 15176 17440 15492 17441
rect 15176 17376 15182 17440
rect 15246 17376 15262 17440
rect 15326 17376 15342 17440
rect 15406 17376 15422 17440
rect 15486 17376 15492 17440
rect 15176 17375 15492 17376
rect 20604 17440 20920 17441
rect 20604 17376 20610 17440
rect 20674 17376 20690 17440
rect 20754 17376 20770 17440
rect 20834 17376 20850 17440
rect 20914 17376 20920 17440
rect 20604 17375 20920 17376
rect 3660 16896 3976 16897
rect 3660 16832 3666 16896
rect 3730 16832 3746 16896
rect 3810 16832 3826 16896
rect 3890 16832 3906 16896
rect 3970 16832 3976 16896
rect 3660 16831 3976 16832
rect 9088 16896 9404 16897
rect 9088 16832 9094 16896
rect 9158 16832 9174 16896
rect 9238 16832 9254 16896
rect 9318 16832 9334 16896
rect 9398 16832 9404 16896
rect 9088 16831 9404 16832
rect 14516 16896 14832 16897
rect 14516 16832 14522 16896
rect 14586 16832 14602 16896
rect 14666 16832 14682 16896
rect 14746 16832 14762 16896
rect 14826 16832 14832 16896
rect 14516 16831 14832 16832
rect 19944 16896 20260 16897
rect 19944 16832 19950 16896
rect 20014 16832 20030 16896
rect 20094 16832 20110 16896
rect 20174 16832 20190 16896
rect 20254 16832 20260 16896
rect 19944 16831 20260 16832
rect 4320 16352 4636 16353
rect 4320 16288 4326 16352
rect 4390 16288 4406 16352
rect 4470 16288 4486 16352
rect 4550 16288 4566 16352
rect 4630 16288 4636 16352
rect 4320 16287 4636 16288
rect 9748 16352 10064 16353
rect 9748 16288 9754 16352
rect 9818 16288 9834 16352
rect 9898 16288 9914 16352
rect 9978 16288 9994 16352
rect 10058 16288 10064 16352
rect 9748 16287 10064 16288
rect 15176 16352 15492 16353
rect 15176 16288 15182 16352
rect 15246 16288 15262 16352
rect 15326 16288 15342 16352
rect 15406 16288 15422 16352
rect 15486 16288 15492 16352
rect 15176 16287 15492 16288
rect 20604 16352 20920 16353
rect 20604 16288 20610 16352
rect 20674 16288 20690 16352
rect 20754 16288 20770 16352
rect 20834 16288 20850 16352
rect 20914 16288 20920 16352
rect 20604 16287 20920 16288
rect 3660 15808 3976 15809
rect 3660 15744 3666 15808
rect 3730 15744 3746 15808
rect 3810 15744 3826 15808
rect 3890 15744 3906 15808
rect 3970 15744 3976 15808
rect 3660 15743 3976 15744
rect 9088 15808 9404 15809
rect 9088 15744 9094 15808
rect 9158 15744 9174 15808
rect 9238 15744 9254 15808
rect 9318 15744 9334 15808
rect 9398 15744 9404 15808
rect 9088 15743 9404 15744
rect 14516 15808 14832 15809
rect 14516 15744 14522 15808
rect 14586 15744 14602 15808
rect 14666 15744 14682 15808
rect 14746 15744 14762 15808
rect 14826 15744 14832 15808
rect 14516 15743 14832 15744
rect 19944 15808 20260 15809
rect 19944 15744 19950 15808
rect 20014 15744 20030 15808
rect 20094 15744 20110 15808
rect 20174 15744 20190 15808
rect 20254 15744 20260 15808
rect 19944 15743 20260 15744
rect 4320 15264 4636 15265
rect 4320 15200 4326 15264
rect 4390 15200 4406 15264
rect 4470 15200 4486 15264
rect 4550 15200 4566 15264
rect 4630 15200 4636 15264
rect 4320 15199 4636 15200
rect 9748 15264 10064 15265
rect 9748 15200 9754 15264
rect 9818 15200 9834 15264
rect 9898 15200 9914 15264
rect 9978 15200 9994 15264
rect 10058 15200 10064 15264
rect 9748 15199 10064 15200
rect 15176 15264 15492 15265
rect 15176 15200 15182 15264
rect 15246 15200 15262 15264
rect 15326 15200 15342 15264
rect 15406 15200 15422 15264
rect 15486 15200 15492 15264
rect 15176 15199 15492 15200
rect 20604 15264 20920 15265
rect 20604 15200 20610 15264
rect 20674 15200 20690 15264
rect 20754 15200 20770 15264
rect 20834 15200 20850 15264
rect 20914 15200 20920 15264
rect 20604 15199 20920 15200
rect 3660 14720 3976 14721
rect 3660 14656 3666 14720
rect 3730 14656 3746 14720
rect 3810 14656 3826 14720
rect 3890 14656 3906 14720
rect 3970 14656 3976 14720
rect 3660 14655 3976 14656
rect 9088 14720 9404 14721
rect 9088 14656 9094 14720
rect 9158 14656 9174 14720
rect 9238 14656 9254 14720
rect 9318 14656 9334 14720
rect 9398 14656 9404 14720
rect 9088 14655 9404 14656
rect 14516 14720 14832 14721
rect 14516 14656 14522 14720
rect 14586 14656 14602 14720
rect 14666 14656 14682 14720
rect 14746 14656 14762 14720
rect 14826 14656 14832 14720
rect 14516 14655 14832 14656
rect 19944 14720 20260 14721
rect 19944 14656 19950 14720
rect 20014 14656 20030 14720
rect 20094 14656 20110 14720
rect 20174 14656 20190 14720
rect 20254 14656 20260 14720
rect 19944 14655 20260 14656
rect 4320 14176 4636 14177
rect 4320 14112 4326 14176
rect 4390 14112 4406 14176
rect 4470 14112 4486 14176
rect 4550 14112 4566 14176
rect 4630 14112 4636 14176
rect 4320 14111 4636 14112
rect 9748 14176 10064 14177
rect 9748 14112 9754 14176
rect 9818 14112 9834 14176
rect 9898 14112 9914 14176
rect 9978 14112 9994 14176
rect 10058 14112 10064 14176
rect 9748 14111 10064 14112
rect 15176 14176 15492 14177
rect 15176 14112 15182 14176
rect 15246 14112 15262 14176
rect 15326 14112 15342 14176
rect 15406 14112 15422 14176
rect 15486 14112 15492 14176
rect 15176 14111 15492 14112
rect 20604 14176 20920 14177
rect 20604 14112 20610 14176
rect 20674 14112 20690 14176
rect 20754 14112 20770 14176
rect 20834 14112 20850 14176
rect 20914 14112 20920 14176
rect 20604 14111 20920 14112
rect 3660 13632 3976 13633
rect 3660 13568 3666 13632
rect 3730 13568 3746 13632
rect 3810 13568 3826 13632
rect 3890 13568 3906 13632
rect 3970 13568 3976 13632
rect 3660 13567 3976 13568
rect 9088 13632 9404 13633
rect 9088 13568 9094 13632
rect 9158 13568 9174 13632
rect 9238 13568 9254 13632
rect 9318 13568 9334 13632
rect 9398 13568 9404 13632
rect 9088 13567 9404 13568
rect 14516 13632 14832 13633
rect 14516 13568 14522 13632
rect 14586 13568 14602 13632
rect 14666 13568 14682 13632
rect 14746 13568 14762 13632
rect 14826 13568 14832 13632
rect 14516 13567 14832 13568
rect 19944 13632 20260 13633
rect 19944 13568 19950 13632
rect 20014 13568 20030 13632
rect 20094 13568 20110 13632
rect 20174 13568 20190 13632
rect 20254 13568 20260 13632
rect 19944 13567 20260 13568
rect 4320 13088 4636 13089
rect 4320 13024 4326 13088
rect 4390 13024 4406 13088
rect 4470 13024 4486 13088
rect 4550 13024 4566 13088
rect 4630 13024 4636 13088
rect 4320 13023 4636 13024
rect 9748 13088 10064 13089
rect 9748 13024 9754 13088
rect 9818 13024 9834 13088
rect 9898 13024 9914 13088
rect 9978 13024 9994 13088
rect 10058 13024 10064 13088
rect 9748 13023 10064 13024
rect 15176 13088 15492 13089
rect 15176 13024 15182 13088
rect 15246 13024 15262 13088
rect 15326 13024 15342 13088
rect 15406 13024 15422 13088
rect 15486 13024 15492 13088
rect 15176 13023 15492 13024
rect 20604 13088 20920 13089
rect 20604 13024 20610 13088
rect 20674 13024 20690 13088
rect 20754 13024 20770 13088
rect 20834 13024 20850 13088
rect 20914 13024 20920 13088
rect 20604 13023 20920 13024
rect 3660 12544 3976 12545
rect 3660 12480 3666 12544
rect 3730 12480 3746 12544
rect 3810 12480 3826 12544
rect 3890 12480 3906 12544
rect 3970 12480 3976 12544
rect 3660 12479 3976 12480
rect 9088 12544 9404 12545
rect 9088 12480 9094 12544
rect 9158 12480 9174 12544
rect 9238 12480 9254 12544
rect 9318 12480 9334 12544
rect 9398 12480 9404 12544
rect 9088 12479 9404 12480
rect 14516 12544 14832 12545
rect 14516 12480 14522 12544
rect 14586 12480 14602 12544
rect 14666 12480 14682 12544
rect 14746 12480 14762 12544
rect 14826 12480 14832 12544
rect 14516 12479 14832 12480
rect 19944 12544 20260 12545
rect 19944 12480 19950 12544
rect 20014 12480 20030 12544
rect 20094 12480 20110 12544
rect 20174 12480 20190 12544
rect 20254 12480 20260 12544
rect 19944 12479 20260 12480
rect 4320 12000 4636 12001
rect 4320 11936 4326 12000
rect 4390 11936 4406 12000
rect 4470 11936 4486 12000
rect 4550 11936 4566 12000
rect 4630 11936 4636 12000
rect 4320 11935 4636 11936
rect 9748 12000 10064 12001
rect 9748 11936 9754 12000
rect 9818 11936 9834 12000
rect 9898 11936 9914 12000
rect 9978 11936 9994 12000
rect 10058 11936 10064 12000
rect 9748 11935 10064 11936
rect 15176 12000 15492 12001
rect 15176 11936 15182 12000
rect 15246 11936 15262 12000
rect 15326 11936 15342 12000
rect 15406 11936 15422 12000
rect 15486 11936 15492 12000
rect 15176 11935 15492 11936
rect 20604 12000 20920 12001
rect 20604 11936 20610 12000
rect 20674 11936 20690 12000
rect 20754 11936 20770 12000
rect 20834 11936 20850 12000
rect 20914 11936 20920 12000
rect 20604 11935 20920 11936
rect 3660 11456 3976 11457
rect 3660 11392 3666 11456
rect 3730 11392 3746 11456
rect 3810 11392 3826 11456
rect 3890 11392 3906 11456
rect 3970 11392 3976 11456
rect 3660 11391 3976 11392
rect 9088 11456 9404 11457
rect 9088 11392 9094 11456
rect 9158 11392 9174 11456
rect 9238 11392 9254 11456
rect 9318 11392 9334 11456
rect 9398 11392 9404 11456
rect 9088 11391 9404 11392
rect 14516 11456 14832 11457
rect 14516 11392 14522 11456
rect 14586 11392 14602 11456
rect 14666 11392 14682 11456
rect 14746 11392 14762 11456
rect 14826 11392 14832 11456
rect 14516 11391 14832 11392
rect 19944 11456 20260 11457
rect 19944 11392 19950 11456
rect 20014 11392 20030 11456
rect 20094 11392 20110 11456
rect 20174 11392 20190 11456
rect 20254 11392 20260 11456
rect 19944 11391 20260 11392
rect 4320 10912 4636 10913
rect 4320 10848 4326 10912
rect 4390 10848 4406 10912
rect 4470 10848 4486 10912
rect 4550 10848 4566 10912
rect 4630 10848 4636 10912
rect 4320 10847 4636 10848
rect 9748 10912 10064 10913
rect 9748 10848 9754 10912
rect 9818 10848 9834 10912
rect 9898 10848 9914 10912
rect 9978 10848 9994 10912
rect 10058 10848 10064 10912
rect 9748 10847 10064 10848
rect 15176 10912 15492 10913
rect 15176 10848 15182 10912
rect 15246 10848 15262 10912
rect 15326 10848 15342 10912
rect 15406 10848 15422 10912
rect 15486 10848 15492 10912
rect 15176 10847 15492 10848
rect 20604 10912 20920 10913
rect 20604 10848 20610 10912
rect 20674 10848 20690 10912
rect 20754 10848 20770 10912
rect 20834 10848 20850 10912
rect 20914 10848 20920 10912
rect 20604 10847 20920 10848
rect 3660 10368 3976 10369
rect 3660 10304 3666 10368
rect 3730 10304 3746 10368
rect 3810 10304 3826 10368
rect 3890 10304 3906 10368
rect 3970 10304 3976 10368
rect 3660 10303 3976 10304
rect 9088 10368 9404 10369
rect 9088 10304 9094 10368
rect 9158 10304 9174 10368
rect 9238 10304 9254 10368
rect 9318 10304 9334 10368
rect 9398 10304 9404 10368
rect 9088 10303 9404 10304
rect 14516 10368 14832 10369
rect 14516 10304 14522 10368
rect 14586 10304 14602 10368
rect 14666 10304 14682 10368
rect 14746 10304 14762 10368
rect 14826 10304 14832 10368
rect 14516 10303 14832 10304
rect 19944 10368 20260 10369
rect 19944 10304 19950 10368
rect 20014 10304 20030 10368
rect 20094 10304 20110 10368
rect 20174 10304 20190 10368
rect 20254 10304 20260 10368
rect 19944 10303 20260 10304
rect 22369 10298 22435 10301
rect 23200 10298 24000 10328
rect 22369 10296 24000 10298
rect 22369 10240 22374 10296
rect 22430 10240 24000 10296
rect 22369 10238 24000 10240
rect 22369 10235 22435 10238
rect 23200 10208 24000 10238
rect 4320 9824 4636 9825
rect 4320 9760 4326 9824
rect 4390 9760 4406 9824
rect 4470 9760 4486 9824
rect 4550 9760 4566 9824
rect 4630 9760 4636 9824
rect 4320 9759 4636 9760
rect 9748 9824 10064 9825
rect 9748 9760 9754 9824
rect 9818 9760 9834 9824
rect 9898 9760 9914 9824
rect 9978 9760 9994 9824
rect 10058 9760 10064 9824
rect 9748 9759 10064 9760
rect 15176 9824 15492 9825
rect 15176 9760 15182 9824
rect 15246 9760 15262 9824
rect 15326 9760 15342 9824
rect 15406 9760 15422 9824
rect 15486 9760 15492 9824
rect 15176 9759 15492 9760
rect 20604 9824 20920 9825
rect 20604 9760 20610 9824
rect 20674 9760 20690 9824
rect 20754 9760 20770 9824
rect 20834 9760 20850 9824
rect 20914 9760 20920 9824
rect 20604 9759 20920 9760
rect 3660 9280 3976 9281
rect 3660 9216 3666 9280
rect 3730 9216 3746 9280
rect 3810 9216 3826 9280
rect 3890 9216 3906 9280
rect 3970 9216 3976 9280
rect 3660 9215 3976 9216
rect 9088 9280 9404 9281
rect 9088 9216 9094 9280
rect 9158 9216 9174 9280
rect 9238 9216 9254 9280
rect 9318 9216 9334 9280
rect 9398 9216 9404 9280
rect 9088 9215 9404 9216
rect 14516 9280 14832 9281
rect 14516 9216 14522 9280
rect 14586 9216 14602 9280
rect 14666 9216 14682 9280
rect 14746 9216 14762 9280
rect 14826 9216 14832 9280
rect 14516 9215 14832 9216
rect 19944 9280 20260 9281
rect 19944 9216 19950 9280
rect 20014 9216 20030 9280
rect 20094 9216 20110 9280
rect 20174 9216 20190 9280
rect 20254 9216 20260 9280
rect 19944 9215 20260 9216
rect 0 8938 800 8968
rect 933 8938 999 8941
rect 0 8936 999 8938
rect 0 8880 938 8936
rect 994 8880 999 8936
rect 0 8878 999 8880
rect 0 8848 800 8878
rect 933 8875 999 8878
rect 4320 8736 4636 8737
rect 4320 8672 4326 8736
rect 4390 8672 4406 8736
rect 4470 8672 4486 8736
rect 4550 8672 4566 8736
rect 4630 8672 4636 8736
rect 4320 8671 4636 8672
rect 9748 8736 10064 8737
rect 9748 8672 9754 8736
rect 9818 8672 9834 8736
rect 9898 8672 9914 8736
rect 9978 8672 9994 8736
rect 10058 8672 10064 8736
rect 9748 8671 10064 8672
rect 15176 8736 15492 8737
rect 15176 8672 15182 8736
rect 15246 8672 15262 8736
rect 15326 8672 15342 8736
rect 15406 8672 15422 8736
rect 15486 8672 15492 8736
rect 15176 8671 15492 8672
rect 20604 8736 20920 8737
rect 20604 8672 20610 8736
rect 20674 8672 20690 8736
rect 20754 8672 20770 8736
rect 20834 8672 20850 8736
rect 20914 8672 20920 8736
rect 20604 8671 20920 8672
rect 3660 8192 3976 8193
rect 3660 8128 3666 8192
rect 3730 8128 3746 8192
rect 3810 8128 3826 8192
rect 3890 8128 3906 8192
rect 3970 8128 3976 8192
rect 3660 8127 3976 8128
rect 9088 8192 9404 8193
rect 9088 8128 9094 8192
rect 9158 8128 9174 8192
rect 9238 8128 9254 8192
rect 9318 8128 9334 8192
rect 9398 8128 9404 8192
rect 9088 8127 9404 8128
rect 14516 8192 14832 8193
rect 14516 8128 14522 8192
rect 14586 8128 14602 8192
rect 14666 8128 14682 8192
rect 14746 8128 14762 8192
rect 14826 8128 14832 8192
rect 14516 8127 14832 8128
rect 19944 8192 20260 8193
rect 19944 8128 19950 8192
rect 20014 8128 20030 8192
rect 20094 8128 20110 8192
rect 20174 8128 20190 8192
rect 20254 8128 20260 8192
rect 19944 8127 20260 8128
rect 4320 7648 4636 7649
rect 4320 7584 4326 7648
rect 4390 7584 4406 7648
rect 4470 7584 4486 7648
rect 4550 7584 4566 7648
rect 4630 7584 4636 7648
rect 4320 7583 4636 7584
rect 9748 7648 10064 7649
rect 9748 7584 9754 7648
rect 9818 7584 9834 7648
rect 9898 7584 9914 7648
rect 9978 7584 9994 7648
rect 10058 7584 10064 7648
rect 9748 7583 10064 7584
rect 15176 7648 15492 7649
rect 15176 7584 15182 7648
rect 15246 7584 15262 7648
rect 15326 7584 15342 7648
rect 15406 7584 15422 7648
rect 15486 7584 15492 7648
rect 15176 7583 15492 7584
rect 20604 7648 20920 7649
rect 20604 7584 20610 7648
rect 20674 7584 20690 7648
rect 20754 7584 20770 7648
rect 20834 7584 20850 7648
rect 20914 7584 20920 7648
rect 20604 7583 20920 7584
rect 3660 7104 3976 7105
rect 3660 7040 3666 7104
rect 3730 7040 3746 7104
rect 3810 7040 3826 7104
rect 3890 7040 3906 7104
rect 3970 7040 3976 7104
rect 3660 7039 3976 7040
rect 9088 7104 9404 7105
rect 9088 7040 9094 7104
rect 9158 7040 9174 7104
rect 9238 7040 9254 7104
rect 9318 7040 9334 7104
rect 9398 7040 9404 7104
rect 9088 7039 9404 7040
rect 14516 7104 14832 7105
rect 14516 7040 14522 7104
rect 14586 7040 14602 7104
rect 14666 7040 14682 7104
rect 14746 7040 14762 7104
rect 14826 7040 14832 7104
rect 14516 7039 14832 7040
rect 19944 7104 20260 7105
rect 19944 7040 19950 7104
rect 20014 7040 20030 7104
rect 20094 7040 20110 7104
rect 20174 7040 20190 7104
rect 20254 7040 20260 7104
rect 19944 7039 20260 7040
rect 4320 6560 4636 6561
rect 4320 6496 4326 6560
rect 4390 6496 4406 6560
rect 4470 6496 4486 6560
rect 4550 6496 4566 6560
rect 4630 6496 4636 6560
rect 4320 6495 4636 6496
rect 9748 6560 10064 6561
rect 9748 6496 9754 6560
rect 9818 6496 9834 6560
rect 9898 6496 9914 6560
rect 9978 6496 9994 6560
rect 10058 6496 10064 6560
rect 9748 6495 10064 6496
rect 15176 6560 15492 6561
rect 15176 6496 15182 6560
rect 15246 6496 15262 6560
rect 15326 6496 15342 6560
rect 15406 6496 15422 6560
rect 15486 6496 15492 6560
rect 15176 6495 15492 6496
rect 20604 6560 20920 6561
rect 20604 6496 20610 6560
rect 20674 6496 20690 6560
rect 20754 6496 20770 6560
rect 20834 6496 20850 6560
rect 20914 6496 20920 6560
rect 20604 6495 20920 6496
rect 3660 6016 3976 6017
rect 3660 5952 3666 6016
rect 3730 5952 3746 6016
rect 3810 5952 3826 6016
rect 3890 5952 3906 6016
rect 3970 5952 3976 6016
rect 3660 5951 3976 5952
rect 9088 6016 9404 6017
rect 9088 5952 9094 6016
rect 9158 5952 9174 6016
rect 9238 5952 9254 6016
rect 9318 5952 9334 6016
rect 9398 5952 9404 6016
rect 9088 5951 9404 5952
rect 14516 6016 14832 6017
rect 14516 5952 14522 6016
rect 14586 5952 14602 6016
rect 14666 5952 14682 6016
rect 14746 5952 14762 6016
rect 14826 5952 14832 6016
rect 14516 5951 14832 5952
rect 19944 6016 20260 6017
rect 19944 5952 19950 6016
rect 20014 5952 20030 6016
rect 20094 5952 20110 6016
rect 20174 5952 20190 6016
rect 20254 5952 20260 6016
rect 19944 5951 20260 5952
rect 4320 5472 4636 5473
rect 4320 5408 4326 5472
rect 4390 5408 4406 5472
rect 4470 5408 4486 5472
rect 4550 5408 4566 5472
rect 4630 5408 4636 5472
rect 4320 5407 4636 5408
rect 9748 5472 10064 5473
rect 9748 5408 9754 5472
rect 9818 5408 9834 5472
rect 9898 5408 9914 5472
rect 9978 5408 9994 5472
rect 10058 5408 10064 5472
rect 9748 5407 10064 5408
rect 15176 5472 15492 5473
rect 15176 5408 15182 5472
rect 15246 5408 15262 5472
rect 15326 5408 15342 5472
rect 15406 5408 15422 5472
rect 15486 5408 15492 5472
rect 15176 5407 15492 5408
rect 20604 5472 20920 5473
rect 20604 5408 20610 5472
rect 20674 5408 20690 5472
rect 20754 5408 20770 5472
rect 20834 5408 20850 5472
rect 20914 5408 20920 5472
rect 20604 5407 20920 5408
rect 3660 4928 3976 4929
rect 3660 4864 3666 4928
rect 3730 4864 3746 4928
rect 3810 4864 3826 4928
rect 3890 4864 3906 4928
rect 3970 4864 3976 4928
rect 3660 4863 3976 4864
rect 9088 4928 9404 4929
rect 9088 4864 9094 4928
rect 9158 4864 9174 4928
rect 9238 4864 9254 4928
rect 9318 4864 9334 4928
rect 9398 4864 9404 4928
rect 9088 4863 9404 4864
rect 14516 4928 14832 4929
rect 14516 4864 14522 4928
rect 14586 4864 14602 4928
rect 14666 4864 14682 4928
rect 14746 4864 14762 4928
rect 14826 4864 14832 4928
rect 14516 4863 14832 4864
rect 19944 4928 20260 4929
rect 19944 4864 19950 4928
rect 20014 4864 20030 4928
rect 20094 4864 20110 4928
rect 20174 4864 20190 4928
rect 20254 4864 20260 4928
rect 19944 4863 20260 4864
rect 4320 4384 4636 4385
rect 4320 4320 4326 4384
rect 4390 4320 4406 4384
rect 4470 4320 4486 4384
rect 4550 4320 4566 4384
rect 4630 4320 4636 4384
rect 4320 4319 4636 4320
rect 9748 4384 10064 4385
rect 9748 4320 9754 4384
rect 9818 4320 9834 4384
rect 9898 4320 9914 4384
rect 9978 4320 9994 4384
rect 10058 4320 10064 4384
rect 9748 4319 10064 4320
rect 15176 4384 15492 4385
rect 15176 4320 15182 4384
rect 15246 4320 15262 4384
rect 15326 4320 15342 4384
rect 15406 4320 15422 4384
rect 15486 4320 15492 4384
rect 15176 4319 15492 4320
rect 20604 4384 20920 4385
rect 20604 4320 20610 4384
rect 20674 4320 20690 4384
rect 20754 4320 20770 4384
rect 20834 4320 20850 4384
rect 20914 4320 20920 4384
rect 20604 4319 20920 4320
rect 3660 3840 3976 3841
rect 3660 3776 3666 3840
rect 3730 3776 3746 3840
rect 3810 3776 3826 3840
rect 3890 3776 3906 3840
rect 3970 3776 3976 3840
rect 3660 3775 3976 3776
rect 9088 3840 9404 3841
rect 9088 3776 9094 3840
rect 9158 3776 9174 3840
rect 9238 3776 9254 3840
rect 9318 3776 9334 3840
rect 9398 3776 9404 3840
rect 9088 3775 9404 3776
rect 14516 3840 14832 3841
rect 14516 3776 14522 3840
rect 14586 3776 14602 3840
rect 14666 3776 14682 3840
rect 14746 3776 14762 3840
rect 14826 3776 14832 3840
rect 14516 3775 14832 3776
rect 19944 3840 20260 3841
rect 19944 3776 19950 3840
rect 20014 3776 20030 3840
rect 20094 3776 20110 3840
rect 20174 3776 20190 3840
rect 20254 3776 20260 3840
rect 19944 3775 20260 3776
rect 4320 3296 4636 3297
rect 4320 3232 4326 3296
rect 4390 3232 4406 3296
rect 4470 3232 4486 3296
rect 4550 3232 4566 3296
rect 4630 3232 4636 3296
rect 4320 3231 4636 3232
rect 9748 3296 10064 3297
rect 9748 3232 9754 3296
rect 9818 3232 9834 3296
rect 9898 3232 9914 3296
rect 9978 3232 9994 3296
rect 10058 3232 10064 3296
rect 9748 3231 10064 3232
rect 15176 3296 15492 3297
rect 15176 3232 15182 3296
rect 15246 3232 15262 3296
rect 15326 3232 15342 3296
rect 15406 3232 15422 3296
rect 15486 3232 15492 3296
rect 15176 3231 15492 3232
rect 20604 3296 20920 3297
rect 20604 3232 20610 3296
rect 20674 3232 20690 3296
rect 20754 3232 20770 3296
rect 20834 3232 20850 3296
rect 20914 3232 20920 3296
rect 20604 3231 20920 3232
rect 3660 2752 3976 2753
rect 3660 2688 3666 2752
rect 3730 2688 3746 2752
rect 3810 2688 3826 2752
rect 3890 2688 3906 2752
rect 3970 2688 3976 2752
rect 3660 2687 3976 2688
rect 9088 2752 9404 2753
rect 9088 2688 9094 2752
rect 9158 2688 9174 2752
rect 9238 2688 9254 2752
rect 9318 2688 9334 2752
rect 9398 2688 9404 2752
rect 9088 2687 9404 2688
rect 14516 2752 14832 2753
rect 14516 2688 14522 2752
rect 14586 2688 14602 2752
rect 14666 2688 14682 2752
rect 14746 2688 14762 2752
rect 14826 2688 14832 2752
rect 14516 2687 14832 2688
rect 19944 2752 20260 2753
rect 19944 2688 19950 2752
rect 20014 2688 20030 2752
rect 20094 2688 20110 2752
rect 20174 2688 20190 2752
rect 20254 2688 20260 2752
rect 19944 2687 20260 2688
rect 4320 2208 4636 2209
rect 4320 2144 4326 2208
rect 4390 2144 4406 2208
rect 4470 2144 4486 2208
rect 4550 2144 4566 2208
rect 4630 2144 4636 2208
rect 4320 2143 4636 2144
rect 9748 2208 10064 2209
rect 9748 2144 9754 2208
rect 9818 2144 9834 2208
rect 9898 2144 9914 2208
rect 9978 2144 9994 2208
rect 10058 2144 10064 2208
rect 9748 2143 10064 2144
rect 15176 2208 15492 2209
rect 15176 2144 15182 2208
rect 15246 2144 15262 2208
rect 15326 2144 15342 2208
rect 15406 2144 15422 2208
rect 15486 2144 15492 2208
rect 15176 2143 15492 2144
rect 20604 2208 20920 2209
rect 20604 2144 20610 2208
rect 20674 2144 20690 2208
rect 20754 2144 20770 2208
rect 20834 2144 20850 2208
rect 20914 2144 20920 2208
rect 20604 2143 20920 2144
rect 22829 1458 22895 1461
rect 23200 1458 24000 1488
rect 22829 1456 24000 1458
rect 22829 1400 22834 1456
rect 22890 1400 24000 1456
rect 22829 1398 24000 1400
rect 22829 1395 22895 1398
rect 23200 1368 24000 1398
<< via3 >>
rect 4326 21788 4390 21792
rect 4326 21732 4330 21788
rect 4330 21732 4386 21788
rect 4386 21732 4390 21788
rect 4326 21728 4390 21732
rect 4406 21788 4470 21792
rect 4406 21732 4410 21788
rect 4410 21732 4466 21788
rect 4466 21732 4470 21788
rect 4406 21728 4470 21732
rect 4486 21788 4550 21792
rect 4486 21732 4490 21788
rect 4490 21732 4546 21788
rect 4546 21732 4550 21788
rect 4486 21728 4550 21732
rect 4566 21788 4630 21792
rect 4566 21732 4570 21788
rect 4570 21732 4626 21788
rect 4626 21732 4630 21788
rect 4566 21728 4630 21732
rect 9754 21788 9818 21792
rect 9754 21732 9758 21788
rect 9758 21732 9814 21788
rect 9814 21732 9818 21788
rect 9754 21728 9818 21732
rect 9834 21788 9898 21792
rect 9834 21732 9838 21788
rect 9838 21732 9894 21788
rect 9894 21732 9898 21788
rect 9834 21728 9898 21732
rect 9914 21788 9978 21792
rect 9914 21732 9918 21788
rect 9918 21732 9974 21788
rect 9974 21732 9978 21788
rect 9914 21728 9978 21732
rect 9994 21788 10058 21792
rect 9994 21732 9998 21788
rect 9998 21732 10054 21788
rect 10054 21732 10058 21788
rect 9994 21728 10058 21732
rect 15182 21788 15246 21792
rect 15182 21732 15186 21788
rect 15186 21732 15242 21788
rect 15242 21732 15246 21788
rect 15182 21728 15246 21732
rect 15262 21788 15326 21792
rect 15262 21732 15266 21788
rect 15266 21732 15322 21788
rect 15322 21732 15326 21788
rect 15262 21728 15326 21732
rect 15342 21788 15406 21792
rect 15342 21732 15346 21788
rect 15346 21732 15402 21788
rect 15402 21732 15406 21788
rect 15342 21728 15406 21732
rect 15422 21788 15486 21792
rect 15422 21732 15426 21788
rect 15426 21732 15482 21788
rect 15482 21732 15486 21788
rect 15422 21728 15486 21732
rect 20610 21788 20674 21792
rect 20610 21732 20614 21788
rect 20614 21732 20670 21788
rect 20670 21732 20674 21788
rect 20610 21728 20674 21732
rect 20690 21788 20754 21792
rect 20690 21732 20694 21788
rect 20694 21732 20750 21788
rect 20750 21732 20754 21788
rect 20690 21728 20754 21732
rect 20770 21788 20834 21792
rect 20770 21732 20774 21788
rect 20774 21732 20830 21788
rect 20830 21732 20834 21788
rect 20770 21728 20834 21732
rect 20850 21788 20914 21792
rect 20850 21732 20854 21788
rect 20854 21732 20910 21788
rect 20910 21732 20914 21788
rect 20850 21728 20914 21732
rect 3666 21244 3730 21248
rect 3666 21188 3670 21244
rect 3670 21188 3726 21244
rect 3726 21188 3730 21244
rect 3666 21184 3730 21188
rect 3746 21244 3810 21248
rect 3746 21188 3750 21244
rect 3750 21188 3806 21244
rect 3806 21188 3810 21244
rect 3746 21184 3810 21188
rect 3826 21244 3890 21248
rect 3826 21188 3830 21244
rect 3830 21188 3886 21244
rect 3886 21188 3890 21244
rect 3826 21184 3890 21188
rect 3906 21244 3970 21248
rect 3906 21188 3910 21244
rect 3910 21188 3966 21244
rect 3966 21188 3970 21244
rect 3906 21184 3970 21188
rect 9094 21244 9158 21248
rect 9094 21188 9098 21244
rect 9098 21188 9154 21244
rect 9154 21188 9158 21244
rect 9094 21184 9158 21188
rect 9174 21244 9238 21248
rect 9174 21188 9178 21244
rect 9178 21188 9234 21244
rect 9234 21188 9238 21244
rect 9174 21184 9238 21188
rect 9254 21244 9318 21248
rect 9254 21188 9258 21244
rect 9258 21188 9314 21244
rect 9314 21188 9318 21244
rect 9254 21184 9318 21188
rect 9334 21244 9398 21248
rect 9334 21188 9338 21244
rect 9338 21188 9394 21244
rect 9394 21188 9398 21244
rect 9334 21184 9398 21188
rect 14522 21244 14586 21248
rect 14522 21188 14526 21244
rect 14526 21188 14582 21244
rect 14582 21188 14586 21244
rect 14522 21184 14586 21188
rect 14602 21244 14666 21248
rect 14602 21188 14606 21244
rect 14606 21188 14662 21244
rect 14662 21188 14666 21244
rect 14602 21184 14666 21188
rect 14682 21244 14746 21248
rect 14682 21188 14686 21244
rect 14686 21188 14742 21244
rect 14742 21188 14746 21244
rect 14682 21184 14746 21188
rect 14762 21244 14826 21248
rect 14762 21188 14766 21244
rect 14766 21188 14822 21244
rect 14822 21188 14826 21244
rect 14762 21184 14826 21188
rect 19950 21244 20014 21248
rect 19950 21188 19954 21244
rect 19954 21188 20010 21244
rect 20010 21188 20014 21244
rect 19950 21184 20014 21188
rect 20030 21244 20094 21248
rect 20030 21188 20034 21244
rect 20034 21188 20090 21244
rect 20090 21188 20094 21244
rect 20030 21184 20094 21188
rect 20110 21244 20174 21248
rect 20110 21188 20114 21244
rect 20114 21188 20170 21244
rect 20170 21188 20174 21244
rect 20110 21184 20174 21188
rect 20190 21244 20254 21248
rect 20190 21188 20194 21244
rect 20194 21188 20250 21244
rect 20250 21188 20254 21244
rect 20190 21184 20254 21188
rect 4326 20700 4390 20704
rect 4326 20644 4330 20700
rect 4330 20644 4386 20700
rect 4386 20644 4390 20700
rect 4326 20640 4390 20644
rect 4406 20700 4470 20704
rect 4406 20644 4410 20700
rect 4410 20644 4466 20700
rect 4466 20644 4470 20700
rect 4406 20640 4470 20644
rect 4486 20700 4550 20704
rect 4486 20644 4490 20700
rect 4490 20644 4546 20700
rect 4546 20644 4550 20700
rect 4486 20640 4550 20644
rect 4566 20700 4630 20704
rect 4566 20644 4570 20700
rect 4570 20644 4626 20700
rect 4626 20644 4630 20700
rect 4566 20640 4630 20644
rect 9754 20700 9818 20704
rect 9754 20644 9758 20700
rect 9758 20644 9814 20700
rect 9814 20644 9818 20700
rect 9754 20640 9818 20644
rect 9834 20700 9898 20704
rect 9834 20644 9838 20700
rect 9838 20644 9894 20700
rect 9894 20644 9898 20700
rect 9834 20640 9898 20644
rect 9914 20700 9978 20704
rect 9914 20644 9918 20700
rect 9918 20644 9974 20700
rect 9974 20644 9978 20700
rect 9914 20640 9978 20644
rect 9994 20700 10058 20704
rect 9994 20644 9998 20700
rect 9998 20644 10054 20700
rect 10054 20644 10058 20700
rect 9994 20640 10058 20644
rect 15182 20700 15246 20704
rect 15182 20644 15186 20700
rect 15186 20644 15242 20700
rect 15242 20644 15246 20700
rect 15182 20640 15246 20644
rect 15262 20700 15326 20704
rect 15262 20644 15266 20700
rect 15266 20644 15322 20700
rect 15322 20644 15326 20700
rect 15262 20640 15326 20644
rect 15342 20700 15406 20704
rect 15342 20644 15346 20700
rect 15346 20644 15402 20700
rect 15402 20644 15406 20700
rect 15342 20640 15406 20644
rect 15422 20700 15486 20704
rect 15422 20644 15426 20700
rect 15426 20644 15482 20700
rect 15482 20644 15486 20700
rect 15422 20640 15486 20644
rect 20610 20700 20674 20704
rect 20610 20644 20614 20700
rect 20614 20644 20670 20700
rect 20670 20644 20674 20700
rect 20610 20640 20674 20644
rect 20690 20700 20754 20704
rect 20690 20644 20694 20700
rect 20694 20644 20750 20700
rect 20750 20644 20754 20700
rect 20690 20640 20754 20644
rect 20770 20700 20834 20704
rect 20770 20644 20774 20700
rect 20774 20644 20830 20700
rect 20830 20644 20834 20700
rect 20770 20640 20834 20644
rect 20850 20700 20914 20704
rect 20850 20644 20854 20700
rect 20854 20644 20910 20700
rect 20910 20644 20914 20700
rect 20850 20640 20914 20644
rect 3666 20156 3730 20160
rect 3666 20100 3670 20156
rect 3670 20100 3726 20156
rect 3726 20100 3730 20156
rect 3666 20096 3730 20100
rect 3746 20156 3810 20160
rect 3746 20100 3750 20156
rect 3750 20100 3806 20156
rect 3806 20100 3810 20156
rect 3746 20096 3810 20100
rect 3826 20156 3890 20160
rect 3826 20100 3830 20156
rect 3830 20100 3886 20156
rect 3886 20100 3890 20156
rect 3826 20096 3890 20100
rect 3906 20156 3970 20160
rect 3906 20100 3910 20156
rect 3910 20100 3966 20156
rect 3966 20100 3970 20156
rect 3906 20096 3970 20100
rect 9094 20156 9158 20160
rect 9094 20100 9098 20156
rect 9098 20100 9154 20156
rect 9154 20100 9158 20156
rect 9094 20096 9158 20100
rect 9174 20156 9238 20160
rect 9174 20100 9178 20156
rect 9178 20100 9234 20156
rect 9234 20100 9238 20156
rect 9174 20096 9238 20100
rect 9254 20156 9318 20160
rect 9254 20100 9258 20156
rect 9258 20100 9314 20156
rect 9314 20100 9318 20156
rect 9254 20096 9318 20100
rect 9334 20156 9398 20160
rect 9334 20100 9338 20156
rect 9338 20100 9394 20156
rect 9394 20100 9398 20156
rect 9334 20096 9398 20100
rect 14522 20156 14586 20160
rect 14522 20100 14526 20156
rect 14526 20100 14582 20156
rect 14582 20100 14586 20156
rect 14522 20096 14586 20100
rect 14602 20156 14666 20160
rect 14602 20100 14606 20156
rect 14606 20100 14662 20156
rect 14662 20100 14666 20156
rect 14602 20096 14666 20100
rect 14682 20156 14746 20160
rect 14682 20100 14686 20156
rect 14686 20100 14742 20156
rect 14742 20100 14746 20156
rect 14682 20096 14746 20100
rect 14762 20156 14826 20160
rect 14762 20100 14766 20156
rect 14766 20100 14822 20156
rect 14822 20100 14826 20156
rect 14762 20096 14826 20100
rect 19950 20156 20014 20160
rect 19950 20100 19954 20156
rect 19954 20100 20010 20156
rect 20010 20100 20014 20156
rect 19950 20096 20014 20100
rect 20030 20156 20094 20160
rect 20030 20100 20034 20156
rect 20034 20100 20090 20156
rect 20090 20100 20094 20156
rect 20030 20096 20094 20100
rect 20110 20156 20174 20160
rect 20110 20100 20114 20156
rect 20114 20100 20170 20156
rect 20170 20100 20174 20156
rect 20110 20096 20174 20100
rect 20190 20156 20254 20160
rect 20190 20100 20194 20156
rect 20194 20100 20250 20156
rect 20250 20100 20254 20156
rect 20190 20096 20254 20100
rect 4326 19612 4390 19616
rect 4326 19556 4330 19612
rect 4330 19556 4386 19612
rect 4386 19556 4390 19612
rect 4326 19552 4390 19556
rect 4406 19612 4470 19616
rect 4406 19556 4410 19612
rect 4410 19556 4466 19612
rect 4466 19556 4470 19612
rect 4406 19552 4470 19556
rect 4486 19612 4550 19616
rect 4486 19556 4490 19612
rect 4490 19556 4546 19612
rect 4546 19556 4550 19612
rect 4486 19552 4550 19556
rect 4566 19612 4630 19616
rect 4566 19556 4570 19612
rect 4570 19556 4626 19612
rect 4626 19556 4630 19612
rect 4566 19552 4630 19556
rect 9754 19612 9818 19616
rect 9754 19556 9758 19612
rect 9758 19556 9814 19612
rect 9814 19556 9818 19612
rect 9754 19552 9818 19556
rect 9834 19612 9898 19616
rect 9834 19556 9838 19612
rect 9838 19556 9894 19612
rect 9894 19556 9898 19612
rect 9834 19552 9898 19556
rect 9914 19612 9978 19616
rect 9914 19556 9918 19612
rect 9918 19556 9974 19612
rect 9974 19556 9978 19612
rect 9914 19552 9978 19556
rect 9994 19612 10058 19616
rect 9994 19556 9998 19612
rect 9998 19556 10054 19612
rect 10054 19556 10058 19612
rect 9994 19552 10058 19556
rect 15182 19612 15246 19616
rect 15182 19556 15186 19612
rect 15186 19556 15242 19612
rect 15242 19556 15246 19612
rect 15182 19552 15246 19556
rect 15262 19612 15326 19616
rect 15262 19556 15266 19612
rect 15266 19556 15322 19612
rect 15322 19556 15326 19612
rect 15262 19552 15326 19556
rect 15342 19612 15406 19616
rect 15342 19556 15346 19612
rect 15346 19556 15402 19612
rect 15402 19556 15406 19612
rect 15342 19552 15406 19556
rect 15422 19612 15486 19616
rect 15422 19556 15426 19612
rect 15426 19556 15482 19612
rect 15482 19556 15486 19612
rect 15422 19552 15486 19556
rect 20610 19612 20674 19616
rect 20610 19556 20614 19612
rect 20614 19556 20670 19612
rect 20670 19556 20674 19612
rect 20610 19552 20674 19556
rect 20690 19612 20754 19616
rect 20690 19556 20694 19612
rect 20694 19556 20750 19612
rect 20750 19556 20754 19612
rect 20690 19552 20754 19556
rect 20770 19612 20834 19616
rect 20770 19556 20774 19612
rect 20774 19556 20830 19612
rect 20830 19556 20834 19612
rect 20770 19552 20834 19556
rect 20850 19612 20914 19616
rect 20850 19556 20854 19612
rect 20854 19556 20910 19612
rect 20910 19556 20914 19612
rect 20850 19552 20914 19556
rect 3666 19068 3730 19072
rect 3666 19012 3670 19068
rect 3670 19012 3726 19068
rect 3726 19012 3730 19068
rect 3666 19008 3730 19012
rect 3746 19068 3810 19072
rect 3746 19012 3750 19068
rect 3750 19012 3806 19068
rect 3806 19012 3810 19068
rect 3746 19008 3810 19012
rect 3826 19068 3890 19072
rect 3826 19012 3830 19068
rect 3830 19012 3886 19068
rect 3886 19012 3890 19068
rect 3826 19008 3890 19012
rect 3906 19068 3970 19072
rect 3906 19012 3910 19068
rect 3910 19012 3966 19068
rect 3966 19012 3970 19068
rect 3906 19008 3970 19012
rect 9094 19068 9158 19072
rect 9094 19012 9098 19068
rect 9098 19012 9154 19068
rect 9154 19012 9158 19068
rect 9094 19008 9158 19012
rect 9174 19068 9238 19072
rect 9174 19012 9178 19068
rect 9178 19012 9234 19068
rect 9234 19012 9238 19068
rect 9174 19008 9238 19012
rect 9254 19068 9318 19072
rect 9254 19012 9258 19068
rect 9258 19012 9314 19068
rect 9314 19012 9318 19068
rect 9254 19008 9318 19012
rect 9334 19068 9398 19072
rect 9334 19012 9338 19068
rect 9338 19012 9394 19068
rect 9394 19012 9398 19068
rect 9334 19008 9398 19012
rect 14522 19068 14586 19072
rect 14522 19012 14526 19068
rect 14526 19012 14582 19068
rect 14582 19012 14586 19068
rect 14522 19008 14586 19012
rect 14602 19068 14666 19072
rect 14602 19012 14606 19068
rect 14606 19012 14662 19068
rect 14662 19012 14666 19068
rect 14602 19008 14666 19012
rect 14682 19068 14746 19072
rect 14682 19012 14686 19068
rect 14686 19012 14742 19068
rect 14742 19012 14746 19068
rect 14682 19008 14746 19012
rect 14762 19068 14826 19072
rect 14762 19012 14766 19068
rect 14766 19012 14822 19068
rect 14822 19012 14826 19068
rect 14762 19008 14826 19012
rect 19950 19068 20014 19072
rect 19950 19012 19954 19068
rect 19954 19012 20010 19068
rect 20010 19012 20014 19068
rect 19950 19008 20014 19012
rect 20030 19068 20094 19072
rect 20030 19012 20034 19068
rect 20034 19012 20090 19068
rect 20090 19012 20094 19068
rect 20030 19008 20094 19012
rect 20110 19068 20174 19072
rect 20110 19012 20114 19068
rect 20114 19012 20170 19068
rect 20170 19012 20174 19068
rect 20110 19008 20174 19012
rect 20190 19068 20254 19072
rect 20190 19012 20194 19068
rect 20194 19012 20250 19068
rect 20250 19012 20254 19068
rect 20190 19008 20254 19012
rect 4326 18524 4390 18528
rect 4326 18468 4330 18524
rect 4330 18468 4386 18524
rect 4386 18468 4390 18524
rect 4326 18464 4390 18468
rect 4406 18524 4470 18528
rect 4406 18468 4410 18524
rect 4410 18468 4466 18524
rect 4466 18468 4470 18524
rect 4406 18464 4470 18468
rect 4486 18524 4550 18528
rect 4486 18468 4490 18524
rect 4490 18468 4546 18524
rect 4546 18468 4550 18524
rect 4486 18464 4550 18468
rect 4566 18524 4630 18528
rect 4566 18468 4570 18524
rect 4570 18468 4626 18524
rect 4626 18468 4630 18524
rect 4566 18464 4630 18468
rect 9754 18524 9818 18528
rect 9754 18468 9758 18524
rect 9758 18468 9814 18524
rect 9814 18468 9818 18524
rect 9754 18464 9818 18468
rect 9834 18524 9898 18528
rect 9834 18468 9838 18524
rect 9838 18468 9894 18524
rect 9894 18468 9898 18524
rect 9834 18464 9898 18468
rect 9914 18524 9978 18528
rect 9914 18468 9918 18524
rect 9918 18468 9974 18524
rect 9974 18468 9978 18524
rect 9914 18464 9978 18468
rect 9994 18524 10058 18528
rect 9994 18468 9998 18524
rect 9998 18468 10054 18524
rect 10054 18468 10058 18524
rect 9994 18464 10058 18468
rect 15182 18524 15246 18528
rect 15182 18468 15186 18524
rect 15186 18468 15242 18524
rect 15242 18468 15246 18524
rect 15182 18464 15246 18468
rect 15262 18524 15326 18528
rect 15262 18468 15266 18524
rect 15266 18468 15322 18524
rect 15322 18468 15326 18524
rect 15262 18464 15326 18468
rect 15342 18524 15406 18528
rect 15342 18468 15346 18524
rect 15346 18468 15402 18524
rect 15402 18468 15406 18524
rect 15342 18464 15406 18468
rect 15422 18524 15486 18528
rect 15422 18468 15426 18524
rect 15426 18468 15482 18524
rect 15482 18468 15486 18524
rect 15422 18464 15486 18468
rect 20610 18524 20674 18528
rect 20610 18468 20614 18524
rect 20614 18468 20670 18524
rect 20670 18468 20674 18524
rect 20610 18464 20674 18468
rect 20690 18524 20754 18528
rect 20690 18468 20694 18524
rect 20694 18468 20750 18524
rect 20750 18468 20754 18524
rect 20690 18464 20754 18468
rect 20770 18524 20834 18528
rect 20770 18468 20774 18524
rect 20774 18468 20830 18524
rect 20830 18468 20834 18524
rect 20770 18464 20834 18468
rect 20850 18524 20914 18528
rect 20850 18468 20854 18524
rect 20854 18468 20910 18524
rect 20910 18468 20914 18524
rect 20850 18464 20914 18468
rect 3666 17980 3730 17984
rect 3666 17924 3670 17980
rect 3670 17924 3726 17980
rect 3726 17924 3730 17980
rect 3666 17920 3730 17924
rect 3746 17980 3810 17984
rect 3746 17924 3750 17980
rect 3750 17924 3806 17980
rect 3806 17924 3810 17980
rect 3746 17920 3810 17924
rect 3826 17980 3890 17984
rect 3826 17924 3830 17980
rect 3830 17924 3886 17980
rect 3886 17924 3890 17980
rect 3826 17920 3890 17924
rect 3906 17980 3970 17984
rect 3906 17924 3910 17980
rect 3910 17924 3966 17980
rect 3966 17924 3970 17980
rect 3906 17920 3970 17924
rect 9094 17980 9158 17984
rect 9094 17924 9098 17980
rect 9098 17924 9154 17980
rect 9154 17924 9158 17980
rect 9094 17920 9158 17924
rect 9174 17980 9238 17984
rect 9174 17924 9178 17980
rect 9178 17924 9234 17980
rect 9234 17924 9238 17980
rect 9174 17920 9238 17924
rect 9254 17980 9318 17984
rect 9254 17924 9258 17980
rect 9258 17924 9314 17980
rect 9314 17924 9318 17980
rect 9254 17920 9318 17924
rect 9334 17980 9398 17984
rect 9334 17924 9338 17980
rect 9338 17924 9394 17980
rect 9394 17924 9398 17980
rect 9334 17920 9398 17924
rect 14522 17980 14586 17984
rect 14522 17924 14526 17980
rect 14526 17924 14582 17980
rect 14582 17924 14586 17980
rect 14522 17920 14586 17924
rect 14602 17980 14666 17984
rect 14602 17924 14606 17980
rect 14606 17924 14662 17980
rect 14662 17924 14666 17980
rect 14602 17920 14666 17924
rect 14682 17980 14746 17984
rect 14682 17924 14686 17980
rect 14686 17924 14742 17980
rect 14742 17924 14746 17980
rect 14682 17920 14746 17924
rect 14762 17980 14826 17984
rect 14762 17924 14766 17980
rect 14766 17924 14822 17980
rect 14822 17924 14826 17980
rect 14762 17920 14826 17924
rect 19950 17980 20014 17984
rect 19950 17924 19954 17980
rect 19954 17924 20010 17980
rect 20010 17924 20014 17980
rect 19950 17920 20014 17924
rect 20030 17980 20094 17984
rect 20030 17924 20034 17980
rect 20034 17924 20090 17980
rect 20090 17924 20094 17980
rect 20030 17920 20094 17924
rect 20110 17980 20174 17984
rect 20110 17924 20114 17980
rect 20114 17924 20170 17980
rect 20170 17924 20174 17980
rect 20110 17920 20174 17924
rect 20190 17980 20254 17984
rect 20190 17924 20194 17980
rect 20194 17924 20250 17980
rect 20250 17924 20254 17980
rect 20190 17920 20254 17924
rect 4326 17436 4390 17440
rect 4326 17380 4330 17436
rect 4330 17380 4386 17436
rect 4386 17380 4390 17436
rect 4326 17376 4390 17380
rect 4406 17436 4470 17440
rect 4406 17380 4410 17436
rect 4410 17380 4466 17436
rect 4466 17380 4470 17436
rect 4406 17376 4470 17380
rect 4486 17436 4550 17440
rect 4486 17380 4490 17436
rect 4490 17380 4546 17436
rect 4546 17380 4550 17436
rect 4486 17376 4550 17380
rect 4566 17436 4630 17440
rect 4566 17380 4570 17436
rect 4570 17380 4626 17436
rect 4626 17380 4630 17436
rect 4566 17376 4630 17380
rect 9754 17436 9818 17440
rect 9754 17380 9758 17436
rect 9758 17380 9814 17436
rect 9814 17380 9818 17436
rect 9754 17376 9818 17380
rect 9834 17436 9898 17440
rect 9834 17380 9838 17436
rect 9838 17380 9894 17436
rect 9894 17380 9898 17436
rect 9834 17376 9898 17380
rect 9914 17436 9978 17440
rect 9914 17380 9918 17436
rect 9918 17380 9974 17436
rect 9974 17380 9978 17436
rect 9914 17376 9978 17380
rect 9994 17436 10058 17440
rect 9994 17380 9998 17436
rect 9998 17380 10054 17436
rect 10054 17380 10058 17436
rect 9994 17376 10058 17380
rect 15182 17436 15246 17440
rect 15182 17380 15186 17436
rect 15186 17380 15242 17436
rect 15242 17380 15246 17436
rect 15182 17376 15246 17380
rect 15262 17436 15326 17440
rect 15262 17380 15266 17436
rect 15266 17380 15322 17436
rect 15322 17380 15326 17436
rect 15262 17376 15326 17380
rect 15342 17436 15406 17440
rect 15342 17380 15346 17436
rect 15346 17380 15402 17436
rect 15402 17380 15406 17436
rect 15342 17376 15406 17380
rect 15422 17436 15486 17440
rect 15422 17380 15426 17436
rect 15426 17380 15482 17436
rect 15482 17380 15486 17436
rect 15422 17376 15486 17380
rect 20610 17436 20674 17440
rect 20610 17380 20614 17436
rect 20614 17380 20670 17436
rect 20670 17380 20674 17436
rect 20610 17376 20674 17380
rect 20690 17436 20754 17440
rect 20690 17380 20694 17436
rect 20694 17380 20750 17436
rect 20750 17380 20754 17436
rect 20690 17376 20754 17380
rect 20770 17436 20834 17440
rect 20770 17380 20774 17436
rect 20774 17380 20830 17436
rect 20830 17380 20834 17436
rect 20770 17376 20834 17380
rect 20850 17436 20914 17440
rect 20850 17380 20854 17436
rect 20854 17380 20910 17436
rect 20910 17380 20914 17436
rect 20850 17376 20914 17380
rect 3666 16892 3730 16896
rect 3666 16836 3670 16892
rect 3670 16836 3726 16892
rect 3726 16836 3730 16892
rect 3666 16832 3730 16836
rect 3746 16892 3810 16896
rect 3746 16836 3750 16892
rect 3750 16836 3806 16892
rect 3806 16836 3810 16892
rect 3746 16832 3810 16836
rect 3826 16892 3890 16896
rect 3826 16836 3830 16892
rect 3830 16836 3886 16892
rect 3886 16836 3890 16892
rect 3826 16832 3890 16836
rect 3906 16892 3970 16896
rect 3906 16836 3910 16892
rect 3910 16836 3966 16892
rect 3966 16836 3970 16892
rect 3906 16832 3970 16836
rect 9094 16892 9158 16896
rect 9094 16836 9098 16892
rect 9098 16836 9154 16892
rect 9154 16836 9158 16892
rect 9094 16832 9158 16836
rect 9174 16892 9238 16896
rect 9174 16836 9178 16892
rect 9178 16836 9234 16892
rect 9234 16836 9238 16892
rect 9174 16832 9238 16836
rect 9254 16892 9318 16896
rect 9254 16836 9258 16892
rect 9258 16836 9314 16892
rect 9314 16836 9318 16892
rect 9254 16832 9318 16836
rect 9334 16892 9398 16896
rect 9334 16836 9338 16892
rect 9338 16836 9394 16892
rect 9394 16836 9398 16892
rect 9334 16832 9398 16836
rect 14522 16892 14586 16896
rect 14522 16836 14526 16892
rect 14526 16836 14582 16892
rect 14582 16836 14586 16892
rect 14522 16832 14586 16836
rect 14602 16892 14666 16896
rect 14602 16836 14606 16892
rect 14606 16836 14662 16892
rect 14662 16836 14666 16892
rect 14602 16832 14666 16836
rect 14682 16892 14746 16896
rect 14682 16836 14686 16892
rect 14686 16836 14742 16892
rect 14742 16836 14746 16892
rect 14682 16832 14746 16836
rect 14762 16892 14826 16896
rect 14762 16836 14766 16892
rect 14766 16836 14822 16892
rect 14822 16836 14826 16892
rect 14762 16832 14826 16836
rect 19950 16892 20014 16896
rect 19950 16836 19954 16892
rect 19954 16836 20010 16892
rect 20010 16836 20014 16892
rect 19950 16832 20014 16836
rect 20030 16892 20094 16896
rect 20030 16836 20034 16892
rect 20034 16836 20090 16892
rect 20090 16836 20094 16892
rect 20030 16832 20094 16836
rect 20110 16892 20174 16896
rect 20110 16836 20114 16892
rect 20114 16836 20170 16892
rect 20170 16836 20174 16892
rect 20110 16832 20174 16836
rect 20190 16892 20254 16896
rect 20190 16836 20194 16892
rect 20194 16836 20250 16892
rect 20250 16836 20254 16892
rect 20190 16832 20254 16836
rect 4326 16348 4390 16352
rect 4326 16292 4330 16348
rect 4330 16292 4386 16348
rect 4386 16292 4390 16348
rect 4326 16288 4390 16292
rect 4406 16348 4470 16352
rect 4406 16292 4410 16348
rect 4410 16292 4466 16348
rect 4466 16292 4470 16348
rect 4406 16288 4470 16292
rect 4486 16348 4550 16352
rect 4486 16292 4490 16348
rect 4490 16292 4546 16348
rect 4546 16292 4550 16348
rect 4486 16288 4550 16292
rect 4566 16348 4630 16352
rect 4566 16292 4570 16348
rect 4570 16292 4626 16348
rect 4626 16292 4630 16348
rect 4566 16288 4630 16292
rect 9754 16348 9818 16352
rect 9754 16292 9758 16348
rect 9758 16292 9814 16348
rect 9814 16292 9818 16348
rect 9754 16288 9818 16292
rect 9834 16348 9898 16352
rect 9834 16292 9838 16348
rect 9838 16292 9894 16348
rect 9894 16292 9898 16348
rect 9834 16288 9898 16292
rect 9914 16348 9978 16352
rect 9914 16292 9918 16348
rect 9918 16292 9974 16348
rect 9974 16292 9978 16348
rect 9914 16288 9978 16292
rect 9994 16348 10058 16352
rect 9994 16292 9998 16348
rect 9998 16292 10054 16348
rect 10054 16292 10058 16348
rect 9994 16288 10058 16292
rect 15182 16348 15246 16352
rect 15182 16292 15186 16348
rect 15186 16292 15242 16348
rect 15242 16292 15246 16348
rect 15182 16288 15246 16292
rect 15262 16348 15326 16352
rect 15262 16292 15266 16348
rect 15266 16292 15322 16348
rect 15322 16292 15326 16348
rect 15262 16288 15326 16292
rect 15342 16348 15406 16352
rect 15342 16292 15346 16348
rect 15346 16292 15402 16348
rect 15402 16292 15406 16348
rect 15342 16288 15406 16292
rect 15422 16348 15486 16352
rect 15422 16292 15426 16348
rect 15426 16292 15482 16348
rect 15482 16292 15486 16348
rect 15422 16288 15486 16292
rect 20610 16348 20674 16352
rect 20610 16292 20614 16348
rect 20614 16292 20670 16348
rect 20670 16292 20674 16348
rect 20610 16288 20674 16292
rect 20690 16348 20754 16352
rect 20690 16292 20694 16348
rect 20694 16292 20750 16348
rect 20750 16292 20754 16348
rect 20690 16288 20754 16292
rect 20770 16348 20834 16352
rect 20770 16292 20774 16348
rect 20774 16292 20830 16348
rect 20830 16292 20834 16348
rect 20770 16288 20834 16292
rect 20850 16348 20914 16352
rect 20850 16292 20854 16348
rect 20854 16292 20910 16348
rect 20910 16292 20914 16348
rect 20850 16288 20914 16292
rect 3666 15804 3730 15808
rect 3666 15748 3670 15804
rect 3670 15748 3726 15804
rect 3726 15748 3730 15804
rect 3666 15744 3730 15748
rect 3746 15804 3810 15808
rect 3746 15748 3750 15804
rect 3750 15748 3806 15804
rect 3806 15748 3810 15804
rect 3746 15744 3810 15748
rect 3826 15804 3890 15808
rect 3826 15748 3830 15804
rect 3830 15748 3886 15804
rect 3886 15748 3890 15804
rect 3826 15744 3890 15748
rect 3906 15804 3970 15808
rect 3906 15748 3910 15804
rect 3910 15748 3966 15804
rect 3966 15748 3970 15804
rect 3906 15744 3970 15748
rect 9094 15804 9158 15808
rect 9094 15748 9098 15804
rect 9098 15748 9154 15804
rect 9154 15748 9158 15804
rect 9094 15744 9158 15748
rect 9174 15804 9238 15808
rect 9174 15748 9178 15804
rect 9178 15748 9234 15804
rect 9234 15748 9238 15804
rect 9174 15744 9238 15748
rect 9254 15804 9318 15808
rect 9254 15748 9258 15804
rect 9258 15748 9314 15804
rect 9314 15748 9318 15804
rect 9254 15744 9318 15748
rect 9334 15804 9398 15808
rect 9334 15748 9338 15804
rect 9338 15748 9394 15804
rect 9394 15748 9398 15804
rect 9334 15744 9398 15748
rect 14522 15804 14586 15808
rect 14522 15748 14526 15804
rect 14526 15748 14582 15804
rect 14582 15748 14586 15804
rect 14522 15744 14586 15748
rect 14602 15804 14666 15808
rect 14602 15748 14606 15804
rect 14606 15748 14662 15804
rect 14662 15748 14666 15804
rect 14602 15744 14666 15748
rect 14682 15804 14746 15808
rect 14682 15748 14686 15804
rect 14686 15748 14742 15804
rect 14742 15748 14746 15804
rect 14682 15744 14746 15748
rect 14762 15804 14826 15808
rect 14762 15748 14766 15804
rect 14766 15748 14822 15804
rect 14822 15748 14826 15804
rect 14762 15744 14826 15748
rect 19950 15804 20014 15808
rect 19950 15748 19954 15804
rect 19954 15748 20010 15804
rect 20010 15748 20014 15804
rect 19950 15744 20014 15748
rect 20030 15804 20094 15808
rect 20030 15748 20034 15804
rect 20034 15748 20090 15804
rect 20090 15748 20094 15804
rect 20030 15744 20094 15748
rect 20110 15804 20174 15808
rect 20110 15748 20114 15804
rect 20114 15748 20170 15804
rect 20170 15748 20174 15804
rect 20110 15744 20174 15748
rect 20190 15804 20254 15808
rect 20190 15748 20194 15804
rect 20194 15748 20250 15804
rect 20250 15748 20254 15804
rect 20190 15744 20254 15748
rect 4326 15260 4390 15264
rect 4326 15204 4330 15260
rect 4330 15204 4386 15260
rect 4386 15204 4390 15260
rect 4326 15200 4390 15204
rect 4406 15260 4470 15264
rect 4406 15204 4410 15260
rect 4410 15204 4466 15260
rect 4466 15204 4470 15260
rect 4406 15200 4470 15204
rect 4486 15260 4550 15264
rect 4486 15204 4490 15260
rect 4490 15204 4546 15260
rect 4546 15204 4550 15260
rect 4486 15200 4550 15204
rect 4566 15260 4630 15264
rect 4566 15204 4570 15260
rect 4570 15204 4626 15260
rect 4626 15204 4630 15260
rect 4566 15200 4630 15204
rect 9754 15260 9818 15264
rect 9754 15204 9758 15260
rect 9758 15204 9814 15260
rect 9814 15204 9818 15260
rect 9754 15200 9818 15204
rect 9834 15260 9898 15264
rect 9834 15204 9838 15260
rect 9838 15204 9894 15260
rect 9894 15204 9898 15260
rect 9834 15200 9898 15204
rect 9914 15260 9978 15264
rect 9914 15204 9918 15260
rect 9918 15204 9974 15260
rect 9974 15204 9978 15260
rect 9914 15200 9978 15204
rect 9994 15260 10058 15264
rect 9994 15204 9998 15260
rect 9998 15204 10054 15260
rect 10054 15204 10058 15260
rect 9994 15200 10058 15204
rect 15182 15260 15246 15264
rect 15182 15204 15186 15260
rect 15186 15204 15242 15260
rect 15242 15204 15246 15260
rect 15182 15200 15246 15204
rect 15262 15260 15326 15264
rect 15262 15204 15266 15260
rect 15266 15204 15322 15260
rect 15322 15204 15326 15260
rect 15262 15200 15326 15204
rect 15342 15260 15406 15264
rect 15342 15204 15346 15260
rect 15346 15204 15402 15260
rect 15402 15204 15406 15260
rect 15342 15200 15406 15204
rect 15422 15260 15486 15264
rect 15422 15204 15426 15260
rect 15426 15204 15482 15260
rect 15482 15204 15486 15260
rect 15422 15200 15486 15204
rect 20610 15260 20674 15264
rect 20610 15204 20614 15260
rect 20614 15204 20670 15260
rect 20670 15204 20674 15260
rect 20610 15200 20674 15204
rect 20690 15260 20754 15264
rect 20690 15204 20694 15260
rect 20694 15204 20750 15260
rect 20750 15204 20754 15260
rect 20690 15200 20754 15204
rect 20770 15260 20834 15264
rect 20770 15204 20774 15260
rect 20774 15204 20830 15260
rect 20830 15204 20834 15260
rect 20770 15200 20834 15204
rect 20850 15260 20914 15264
rect 20850 15204 20854 15260
rect 20854 15204 20910 15260
rect 20910 15204 20914 15260
rect 20850 15200 20914 15204
rect 3666 14716 3730 14720
rect 3666 14660 3670 14716
rect 3670 14660 3726 14716
rect 3726 14660 3730 14716
rect 3666 14656 3730 14660
rect 3746 14716 3810 14720
rect 3746 14660 3750 14716
rect 3750 14660 3806 14716
rect 3806 14660 3810 14716
rect 3746 14656 3810 14660
rect 3826 14716 3890 14720
rect 3826 14660 3830 14716
rect 3830 14660 3886 14716
rect 3886 14660 3890 14716
rect 3826 14656 3890 14660
rect 3906 14716 3970 14720
rect 3906 14660 3910 14716
rect 3910 14660 3966 14716
rect 3966 14660 3970 14716
rect 3906 14656 3970 14660
rect 9094 14716 9158 14720
rect 9094 14660 9098 14716
rect 9098 14660 9154 14716
rect 9154 14660 9158 14716
rect 9094 14656 9158 14660
rect 9174 14716 9238 14720
rect 9174 14660 9178 14716
rect 9178 14660 9234 14716
rect 9234 14660 9238 14716
rect 9174 14656 9238 14660
rect 9254 14716 9318 14720
rect 9254 14660 9258 14716
rect 9258 14660 9314 14716
rect 9314 14660 9318 14716
rect 9254 14656 9318 14660
rect 9334 14716 9398 14720
rect 9334 14660 9338 14716
rect 9338 14660 9394 14716
rect 9394 14660 9398 14716
rect 9334 14656 9398 14660
rect 14522 14716 14586 14720
rect 14522 14660 14526 14716
rect 14526 14660 14582 14716
rect 14582 14660 14586 14716
rect 14522 14656 14586 14660
rect 14602 14716 14666 14720
rect 14602 14660 14606 14716
rect 14606 14660 14662 14716
rect 14662 14660 14666 14716
rect 14602 14656 14666 14660
rect 14682 14716 14746 14720
rect 14682 14660 14686 14716
rect 14686 14660 14742 14716
rect 14742 14660 14746 14716
rect 14682 14656 14746 14660
rect 14762 14716 14826 14720
rect 14762 14660 14766 14716
rect 14766 14660 14822 14716
rect 14822 14660 14826 14716
rect 14762 14656 14826 14660
rect 19950 14716 20014 14720
rect 19950 14660 19954 14716
rect 19954 14660 20010 14716
rect 20010 14660 20014 14716
rect 19950 14656 20014 14660
rect 20030 14716 20094 14720
rect 20030 14660 20034 14716
rect 20034 14660 20090 14716
rect 20090 14660 20094 14716
rect 20030 14656 20094 14660
rect 20110 14716 20174 14720
rect 20110 14660 20114 14716
rect 20114 14660 20170 14716
rect 20170 14660 20174 14716
rect 20110 14656 20174 14660
rect 20190 14716 20254 14720
rect 20190 14660 20194 14716
rect 20194 14660 20250 14716
rect 20250 14660 20254 14716
rect 20190 14656 20254 14660
rect 4326 14172 4390 14176
rect 4326 14116 4330 14172
rect 4330 14116 4386 14172
rect 4386 14116 4390 14172
rect 4326 14112 4390 14116
rect 4406 14172 4470 14176
rect 4406 14116 4410 14172
rect 4410 14116 4466 14172
rect 4466 14116 4470 14172
rect 4406 14112 4470 14116
rect 4486 14172 4550 14176
rect 4486 14116 4490 14172
rect 4490 14116 4546 14172
rect 4546 14116 4550 14172
rect 4486 14112 4550 14116
rect 4566 14172 4630 14176
rect 4566 14116 4570 14172
rect 4570 14116 4626 14172
rect 4626 14116 4630 14172
rect 4566 14112 4630 14116
rect 9754 14172 9818 14176
rect 9754 14116 9758 14172
rect 9758 14116 9814 14172
rect 9814 14116 9818 14172
rect 9754 14112 9818 14116
rect 9834 14172 9898 14176
rect 9834 14116 9838 14172
rect 9838 14116 9894 14172
rect 9894 14116 9898 14172
rect 9834 14112 9898 14116
rect 9914 14172 9978 14176
rect 9914 14116 9918 14172
rect 9918 14116 9974 14172
rect 9974 14116 9978 14172
rect 9914 14112 9978 14116
rect 9994 14172 10058 14176
rect 9994 14116 9998 14172
rect 9998 14116 10054 14172
rect 10054 14116 10058 14172
rect 9994 14112 10058 14116
rect 15182 14172 15246 14176
rect 15182 14116 15186 14172
rect 15186 14116 15242 14172
rect 15242 14116 15246 14172
rect 15182 14112 15246 14116
rect 15262 14172 15326 14176
rect 15262 14116 15266 14172
rect 15266 14116 15322 14172
rect 15322 14116 15326 14172
rect 15262 14112 15326 14116
rect 15342 14172 15406 14176
rect 15342 14116 15346 14172
rect 15346 14116 15402 14172
rect 15402 14116 15406 14172
rect 15342 14112 15406 14116
rect 15422 14172 15486 14176
rect 15422 14116 15426 14172
rect 15426 14116 15482 14172
rect 15482 14116 15486 14172
rect 15422 14112 15486 14116
rect 20610 14172 20674 14176
rect 20610 14116 20614 14172
rect 20614 14116 20670 14172
rect 20670 14116 20674 14172
rect 20610 14112 20674 14116
rect 20690 14172 20754 14176
rect 20690 14116 20694 14172
rect 20694 14116 20750 14172
rect 20750 14116 20754 14172
rect 20690 14112 20754 14116
rect 20770 14172 20834 14176
rect 20770 14116 20774 14172
rect 20774 14116 20830 14172
rect 20830 14116 20834 14172
rect 20770 14112 20834 14116
rect 20850 14172 20914 14176
rect 20850 14116 20854 14172
rect 20854 14116 20910 14172
rect 20910 14116 20914 14172
rect 20850 14112 20914 14116
rect 3666 13628 3730 13632
rect 3666 13572 3670 13628
rect 3670 13572 3726 13628
rect 3726 13572 3730 13628
rect 3666 13568 3730 13572
rect 3746 13628 3810 13632
rect 3746 13572 3750 13628
rect 3750 13572 3806 13628
rect 3806 13572 3810 13628
rect 3746 13568 3810 13572
rect 3826 13628 3890 13632
rect 3826 13572 3830 13628
rect 3830 13572 3886 13628
rect 3886 13572 3890 13628
rect 3826 13568 3890 13572
rect 3906 13628 3970 13632
rect 3906 13572 3910 13628
rect 3910 13572 3966 13628
rect 3966 13572 3970 13628
rect 3906 13568 3970 13572
rect 9094 13628 9158 13632
rect 9094 13572 9098 13628
rect 9098 13572 9154 13628
rect 9154 13572 9158 13628
rect 9094 13568 9158 13572
rect 9174 13628 9238 13632
rect 9174 13572 9178 13628
rect 9178 13572 9234 13628
rect 9234 13572 9238 13628
rect 9174 13568 9238 13572
rect 9254 13628 9318 13632
rect 9254 13572 9258 13628
rect 9258 13572 9314 13628
rect 9314 13572 9318 13628
rect 9254 13568 9318 13572
rect 9334 13628 9398 13632
rect 9334 13572 9338 13628
rect 9338 13572 9394 13628
rect 9394 13572 9398 13628
rect 9334 13568 9398 13572
rect 14522 13628 14586 13632
rect 14522 13572 14526 13628
rect 14526 13572 14582 13628
rect 14582 13572 14586 13628
rect 14522 13568 14586 13572
rect 14602 13628 14666 13632
rect 14602 13572 14606 13628
rect 14606 13572 14662 13628
rect 14662 13572 14666 13628
rect 14602 13568 14666 13572
rect 14682 13628 14746 13632
rect 14682 13572 14686 13628
rect 14686 13572 14742 13628
rect 14742 13572 14746 13628
rect 14682 13568 14746 13572
rect 14762 13628 14826 13632
rect 14762 13572 14766 13628
rect 14766 13572 14822 13628
rect 14822 13572 14826 13628
rect 14762 13568 14826 13572
rect 19950 13628 20014 13632
rect 19950 13572 19954 13628
rect 19954 13572 20010 13628
rect 20010 13572 20014 13628
rect 19950 13568 20014 13572
rect 20030 13628 20094 13632
rect 20030 13572 20034 13628
rect 20034 13572 20090 13628
rect 20090 13572 20094 13628
rect 20030 13568 20094 13572
rect 20110 13628 20174 13632
rect 20110 13572 20114 13628
rect 20114 13572 20170 13628
rect 20170 13572 20174 13628
rect 20110 13568 20174 13572
rect 20190 13628 20254 13632
rect 20190 13572 20194 13628
rect 20194 13572 20250 13628
rect 20250 13572 20254 13628
rect 20190 13568 20254 13572
rect 4326 13084 4390 13088
rect 4326 13028 4330 13084
rect 4330 13028 4386 13084
rect 4386 13028 4390 13084
rect 4326 13024 4390 13028
rect 4406 13084 4470 13088
rect 4406 13028 4410 13084
rect 4410 13028 4466 13084
rect 4466 13028 4470 13084
rect 4406 13024 4470 13028
rect 4486 13084 4550 13088
rect 4486 13028 4490 13084
rect 4490 13028 4546 13084
rect 4546 13028 4550 13084
rect 4486 13024 4550 13028
rect 4566 13084 4630 13088
rect 4566 13028 4570 13084
rect 4570 13028 4626 13084
rect 4626 13028 4630 13084
rect 4566 13024 4630 13028
rect 9754 13084 9818 13088
rect 9754 13028 9758 13084
rect 9758 13028 9814 13084
rect 9814 13028 9818 13084
rect 9754 13024 9818 13028
rect 9834 13084 9898 13088
rect 9834 13028 9838 13084
rect 9838 13028 9894 13084
rect 9894 13028 9898 13084
rect 9834 13024 9898 13028
rect 9914 13084 9978 13088
rect 9914 13028 9918 13084
rect 9918 13028 9974 13084
rect 9974 13028 9978 13084
rect 9914 13024 9978 13028
rect 9994 13084 10058 13088
rect 9994 13028 9998 13084
rect 9998 13028 10054 13084
rect 10054 13028 10058 13084
rect 9994 13024 10058 13028
rect 15182 13084 15246 13088
rect 15182 13028 15186 13084
rect 15186 13028 15242 13084
rect 15242 13028 15246 13084
rect 15182 13024 15246 13028
rect 15262 13084 15326 13088
rect 15262 13028 15266 13084
rect 15266 13028 15322 13084
rect 15322 13028 15326 13084
rect 15262 13024 15326 13028
rect 15342 13084 15406 13088
rect 15342 13028 15346 13084
rect 15346 13028 15402 13084
rect 15402 13028 15406 13084
rect 15342 13024 15406 13028
rect 15422 13084 15486 13088
rect 15422 13028 15426 13084
rect 15426 13028 15482 13084
rect 15482 13028 15486 13084
rect 15422 13024 15486 13028
rect 20610 13084 20674 13088
rect 20610 13028 20614 13084
rect 20614 13028 20670 13084
rect 20670 13028 20674 13084
rect 20610 13024 20674 13028
rect 20690 13084 20754 13088
rect 20690 13028 20694 13084
rect 20694 13028 20750 13084
rect 20750 13028 20754 13084
rect 20690 13024 20754 13028
rect 20770 13084 20834 13088
rect 20770 13028 20774 13084
rect 20774 13028 20830 13084
rect 20830 13028 20834 13084
rect 20770 13024 20834 13028
rect 20850 13084 20914 13088
rect 20850 13028 20854 13084
rect 20854 13028 20910 13084
rect 20910 13028 20914 13084
rect 20850 13024 20914 13028
rect 3666 12540 3730 12544
rect 3666 12484 3670 12540
rect 3670 12484 3726 12540
rect 3726 12484 3730 12540
rect 3666 12480 3730 12484
rect 3746 12540 3810 12544
rect 3746 12484 3750 12540
rect 3750 12484 3806 12540
rect 3806 12484 3810 12540
rect 3746 12480 3810 12484
rect 3826 12540 3890 12544
rect 3826 12484 3830 12540
rect 3830 12484 3886 12540
rect 3886 12484 3890 12540
rect 3826 12480 3890 12484
rect 3906 12540 3970 12544
rect 3906 12484 3910 12540
rect 3910 12484 3966 12540
rect 3966 12484 3970 12540
rect 3906 12480 3970 12484
rect 9094 12540 9158 12544
rect 9094 12484 9098 12540
rect 9098 12484 9154 12540
rect 9154 12484 9158 12540
rect 9094 12480 9158 12484
rect 9174 12540 9238 12544
rect 9174 12484 9178 12540
rect 9178 12484 9234 12540
rect 9234 12484 9238 12540
rect 9174 12480 9238 12484
rect 9254 12540 9318 12544
rect 9254 12484 9258 12540
rect 9258 12484 9314 12540
rect 9314 12484 9318 12540
rect 9254 12480 9318 12484
rect 9334 12540 9398 12544
rect 9334 12484 9338 12540
rect 9338 12484 9394 12540
rect 9394 12484 9398 12540
rect 9334 12480 9398 12484
rect 14522 12540 14586 12544
rect 14522 12484 14526 12540
rect 14526 12484 14582 12540
rect 14582 12484 14586 12540
rect 14522 12480 14586 12484
rect 14602 12540 14666 12544
rect 14602 12484 14606 12540
rect 14606 12484 14662 12540
rect 14662 12484 14666 12540
rect 14602 12480 14666 12484
rect 14682 12540 14746 12544
rect 14682 12484 14686 12540
rect 14686 12484 14742 12540
rect 14742 12484 14746 12540
rect 14682 12480 14746 12484
rect 14762 12540 14826 12544
rect 14762 12484 14766 12540
rect 14766 12484 14822 12540
rect 14822 12484 14826 12540
rect 14762 12480 14826 12484
rect 19950 12540 20014 12544
rect 19950 12484 19954 12540
rect 19954 12484 20010 12540
rect 20010 12484 20014 12540
rect 19950 12480 20014 12484
rect 20030 12540 20094 12544
rect 20030 12484 20034 12540
rect 20034 12484 20090 12540
rect 20090 12484 20094 12540
rect 20030 12480 20094 12484
rect 20110 12540 20174 12544
rect 20110 12484 20114 12540
rect 20114 12484 20170 12540
rect 20170 12484 20174 12540
rect 20110 12480 20174 12484
rect 20190 12540 20254 12544
rect 20190 12484 20194 12540
rect 20194 12484 20250 12540
rect 20250 12484 20254 12540
rect 20190 12480 20254 12484
rect 4326 11996 4390 12000
rect 4326 11940 4330 11996
rect 4330 11940 4386 11996
rect 4386 11940 4390 11996
rect 4326 11936 4390 11940
rect 4406 11996 4470 12000
rect 4406 11940 4410 11996
rect 4410 11940 4466 11996
rect 4466 11940 4470 11996
rect 4406 11936 4470 11940
rect 4486 11996 4550 12000
rect 4486 11940 4490 11996
rect 4490 11940 4546 11996
rect 4546 11940 4550 11996
rect 4486 11936 4550 11940
rect 4566 11996 4630 12000
rect 4566 11940 4570 11996
rect 4570 11940 4626 11996
rect 4626 11940 4630 11996
rect 4566 11936 4630 11940
rect 9754 11996 9818 12000
rect 9754 11940 9758 11996
rect 9758 11940 9814 11996
rect 9814 11940 9818 11996
rect 9754 11936 9818 11940
rect 9834 11996 9898 12000
rect 9834 11940 9838 11996
rect 9838 11940 9894 11996
rect 9894 11940 9898 11996
rect 9834 11936 9898 11940
rect 9914 11996 9978 12000
rect 9914 11940 9918 11996
rect 9918 11940 9974 11996
rect 9974 11940 9978 11996
rect 9914 11936 9978 11940
rect 9994 11996 10058 12000
rect 9994 11940 9998 11996
rect 9998 11940 10054 11996
rect 10054 11940 10058 11996
rect 9994 11936 10058 11940
rect 15182 11996 15246 12000
rect 15182 11940 15186 11996
rect 15186 11940 15242 11996
rect 15242 11940 15246 11996
rect 15182 11936 15246 11940
rect 15262 11996 15326 12000
rect 15262 11940 15266 11996
rect 15266 11940 15322 11996
rect 15322 11940 15326 11996
rect 15262 11936 15326 11940
rect 15342 11996 15406 12000
rect 15342 11940 15346 11996
rect 15346 11940 15402 11996
rect 15402 11940 15406 11996
rect 15342 11936 15406 11940
rect 15422 11996 15486 12000
rect 15422 11940 15426 11996
rect 15426 11940 15482 11996
rect 15482 11940 15486 11996
rect 15422 11936 15486 11940
rect 20610 11996 20674 12000
rect 20610 11940 20614 11996
rect 20614 11940 20670 11996
rect 20670 11940 20674 11996
rect 20610 11936 20674 11940
rect 20690 11996 20754 12000
rect 20690 11940 20694 11996
rect 20694 11940 20750 11996
rect 20750 11940 20754 11996
rect 20690 11936 20754 11940
rect 20770 11996 20834 12000
rect 20770 11940 20774 11996
rect 20774 11940 20830 11996
rect 20830 11940 20834 11996
rect 20770 11936 20834 11940
rect 20850 11996 20914 12000
rect 20850 11940 20854 11996
rect 20854 11940 20910 11996
rect 20910 11940 20914 11996
rect 20850 11936 20914 11940
rect 3666 11452 3730 11456
rect 3666 11396 3670 11452
rect 3670 11396 3726 11452
rect 3726 11396 3730 11452
rect 3666 11392 3730 11396
rect 3746 11452 3810 11456
rect 3746 11396 3750 11452
rect 3750 11396 3806 11452
rect 3806 11396 3810 11452
rect 3746 11392 3810 11396
rect 3826 11452 3890 11456
rect 3826 11396 3830 11452
rect 3830 11396 3886 11452
rect 3886 11396 3890 11452
rect 3826 11392 3890 11396
rect 3906 11452 3970 11456
rect 3906 11396 3910 11452
rect 3910 11396 3966 11452
rect 3966 11396 3970 11452
rect 3906 11392 3970 11396
rect 9094 11452 9158 11456
rect 9094 11396 9098 11452
rect 9098 11396 9154 11452
rect 9154 11396 9158 11452
rect 9094 11392 9158 11396
rect 9174 11452 9238 11456
rect 9174 11396 9178 11452
rect 9178 11396 9234 11452
rect 9234 11396 9238 11452
rect 9174 11392 9238 11396
rect 9254 11452 9318 11456
rect 9254 11396 9258 11452
rect 9258 11396 9314 11452
rect 9314 11396 9318 11452
rect 9254 11392 9318 11396
rect 9334 11452 9398 11456
rect 9334 11396 9338 11452
rect 9338 11396 9394 11452
rect 9394 11396 9398 11452
rect 9334 11392 9398 11396
rect 14522 11452 14586 11456
rect 14522 11396 14526 11452
rect 14526 11396 14582 11452
rect 14582 11396 14586 11452
rect 14522 11392 14586 11396
rect 14602 11452 14666 11456
rect 14602 11396 14606 11452
rect 14606 11396 14662 11452
rect 14662 11396 14666 11452
rect 14602 11392 14666 11396
rect 14682 11452 14746 11456
rect 14682 11396 14686 11452
rect 14686 11396 14742 11452
rect 14742 11396 14746 11452
rect 14682 11392 14746 11396
rect 14762 11452 14826 11456
rect 14762 11396 14766 11452
rect 14766 11396 14822 11452
rect 14822 11396 14826 11452
rect 14762 11392 14826 11396
rect 19950 11452 20014 11456
rect 19950 11396 19954 11452
rect 19954 11396 20010 11452
rect 20010 11396 20014 11452
rect 19950 11392 20014 11396
rect 20030 11452 20094 11456
rect 20030 11396 20034 11452
rect 20034 11396 20090 11452
rect 20090 11396 20094 11452
rect 20030 11392 20094 11396
rect 20110 11452 20174 11456
rect 20110 11396 20114 11452
rect 20114 11396 20170 11452
rect 20170 11396 20174 11452
rect 20110 11392 20174 11396
rect 20190 11452 20254 11456
rect 20190 11396 20194 11452
rect 20194 11396 20250 11452
rect 20250 11396 20254 11452
rect 20190 11392 20254 11396
rect 4326 10908 4390 10912
rect 4326 10852 4330 10908
rect 4330 10852 4386 10908
rect 4386 10852 4390 10908
rect 4326 10848 4390 10852
rect 4406 10908 4470 10912
rect 4406 10852 4410 10908
rect 4410 10852 4466 10908
rect 4466 10852 4470 10908
rect 4406 10848 4470 10852
rect 4486 10908 4550 10912
rect 4486 10852 4490 10908
rect 4490 10852 4546 10908
rect 4546 10852 4550 10908
rect 4486 10848 4550 10852
rect 4566 10908 4630 10912
rect 4566 10852 4570 10908
rect 4570 10852 4626 10908
rect 4626 10852 4630 10908
rect 4566 10848 4630 10852
rect 9754 10908 9818 10912
rect 9754 10852 9758 10908
rect 9758 10852 9814 10908
rect 9814 10852 9818 10908
rect 9754 10848 9818 10852
rect 9834 10908 9898 10912
rect 9834 10852 9838 10908
rect 9838 10852 9894 10908
rect 9894 10852 9898 10908
rect 9834 10848 9898 10852
rect 9914 10908 9978 10912
rect 9914 10852 9918 10908
rect 9918 10852 9974 10908
rect 9974 10852 9978 10908
rect 9914 10848 9978 10852
rect 9994 10908 10058 10912
rect 9994 10852 9998 10908
rect 9998 10852 10054 10908
rect 10054 10852 10058 10908
rect 9994 10848 10058 10852
rect 15182 10908 15246 10912
rect 15182 10852 15186 10908
rect 15186 10852 15242 10908
rect 15242 10852 15246 10908
rect 15182 10848 15246 10852
rect 15262 10908 15326 10912
rect 15262 10852 15266 10908
rect 15266 10852 15322 10908
rect 15322 10852 15326 10908
rect 15262 10848 15326 10852
rect 15342 10908 15406 10912
rect 15342 10852 15346 10908
rect 15346 10852 15402 10908
rect 15402 10852 15406 10908
rect 15342 10848 15406 10852
rect 15422 10908 15486 10912
rect 15422 10852 15426 10908
rect 15426 10852 15482 10908
rect 15482 10852 15486 10908
rect 15422 10848 15486 10852
rect 20610 10908 20674 10912
rect 20610 10852 20614 10908
rect 20614 10852 20670 10908
rect 20670 10852 20674 10908
rect 20610 10848 20674 10852
rect 20690 10908 20754 10912
rect 20690 10852 20694 10908
rect 20694 10852 20750 10908
rect 20750 10852 20754 10908
rect 20690 10848 20754 10852
rect 20770 10908 20834 10912
rect 20770 10852 20774 10908
rect 20774 10852 20830 10908
rect 20830 10852 20834 10908
rect 20770 10848 20834 10852
rect 20850 10908 20914 10912
rect 20850 10852 20854 10908
rect 20854 10852 20910 10908
rect 20910 10852 20914 10908
rect 20850 10848 20914 10852
rect 3666 10364 3730 10368
rect 3666 10308 3670 10364
rect 3670 10308 3726 10364
rect 3726 10308 3730 10364
rect 3666 10304 3730 10308
rect 3746 10364 3810 10368
rect 3746 10308 3750 10364
rect 3750 10308 3806 10364
rect 3806 10308 3810 10364
rect 3746 10304 3810 10308
rect 3826 10364 3890 10368
rect 3826 10308 3830 10364
rect 3830 10308 3886 10364
rect 3886 10308 3890 10364
rect 3826 10304 3890 10308
rect 3906 10364 3970 10368
rect 3906 10308 3910 10364
rect 3910 10308 3966 10364
rect 3966 10308 3970 10364
rect 3906 10304 3970 10308
rect 9094 10364 9158 10368
rect 9094 10308 9098 10364
rect 9098 10308 9154 10364
rect 9154 10308 9158 10364
rect 9094 10304 9158 10308
rect 9174 10364 9238 10368
rect 9174 10308 9178 10364
rect 9178 10308 9234 10364
rect 9234 10308 9238 10364
rect 9174 10304 9238 10308
rect 9254 10364 9318 10368
rect 9254 10308 9258 10364
rect 9258 10308 9314 10364
rect 9314 10308 9318 10364
rect 9254 10304 9318 10308
rect 9334 10364 9398 10368
rect 9334 10308 9338 10364
rect 9338 10308 9394 10364
rect 9394 10308 9398 10364
rect 9334 10304 9398 10308
rect 14522 10364 14586 10368
rect 14522 10308 14526 10364
rect 14526 10308 14582 10364
rect 14582 10308 14586 10364
rect 14522 10304 14586 10308
rect 14602 10364 14666 10368
rect 14602 10308 14606 10364
rect 14606 10308 14662 10364
rect 14662 10308 14666 10364
rect 14602 10304 14666 10308
rect 14682 10364 14746 10368
rect 14682 10308 14686 10364
rect 14686 10308 14742 10364
rect 14742 10308 14746 10364
rect 14682 10304 14746 10308
rect 14762 10364 14826 10368
rect 14762 10308 14766 10364
rect 14766 10308 14822 10364
rect 14822 10308 14826 10364
rect 14762 10304 14826 10308
rect 19950 10364 20014 10368
rect 19950 10308 19954 10364
rect 19954 10308 20010 10364
rect 20010 10308 20014 10364
rect 19950 10304 20014 10308
rect 20030 10364 20094 10368
rect 20030 10308 20034 10364
rect 20034 10308 20090 10364
rect 20090 10308 20094 10364
rect 20030 10304 20094 10308
rect 20110 10364 20174 10368
rect 20110 10308 20114 10364
rect 20114 10308 20170 10364
rect 20170 10308 20174 10364
rect 20110 10304 20174 10308
rect 20190 10364 20254 10368
rect 20190 10308 20194 10364
rect 20194 10308 20250 10364
rect 20250 10308 20254 10364
rect 20190 10304 20254 10308
rect 4326 9820 4390 9824
rect 4326 9764 4330 9820
rect 4330 9764 4386 9820
rect 4386 9764 4390 9820
rect 4326 9760 4390 9764
rect 4406 9820 4470 9824
rect 4406 9764 4410 9820
rect 4410 9764 4466 9820
rect 4466 9764 4470 9820
rect 4406 9760 4470 9764
rect 4486 9820 4550 9824
rect 4486 9764 4490 9820
rect 4490 9764 4546 9820
rect 4546 9764 4550 9820
rect 4486 9760 4550 9764
rect 4566 9820 4630 9824
rect 4566 9764 4570 9820
rect 4570 9764 4626 9820
rect 4626 9764 4630 9820
rect 4566 9760 4630 9764
rect 9754 9820 9818 9824
rect 9754 9764 9758 9820
rect 9758 9764 9814 9820
rect 9814 9764 9818 9820
rect 9754 9760 9818 9764
rect 9834 9820 9898 9824
rect 9834 9764 9838 9820
rect 9838 9764 9894 9820
rect 9894 9764 9898 9820
rect 9834 9760 9898 9764
rect 9914 9820 9978 9824
rect 9914 9764 9918 9820
rect 9918 9764 9974 9820
rect 9974 9764 9978 9820
rect 9914 9760 9978 9764
rect 9994 9820 10058 9824
rect 9994 9764 9998 9820
rect 9998 9764 10054 9820
rect 10054 9764 10058 9820
rect 9994 9760 10058 9764
rect 15182 9820 15246 9824
rect 15182 9764 15186 9820
rect 15186 9764 15242 9820
rect 15242 9764 15246 9820
rect 15182 9760 15246 9764
rect 15262 9820 15326 9824
rect 15262 9764 15266 9820
rect 15266 9764 15322 9820
rect 15322 9764 15326 9820
rect 15262 9760 15326 9764
rect 15342 9820 15406 9824
rect 15342 9764 15346 9820
rect 15346 9764 15402 9820
rect 15402 9764 15406 9820
rect 15342 9760 15406 9764
rect 15422 9820 15486 9824
rect 15422 9764 15426 9820
rect 15426 9764 15482 9820
rect 15482 9764 15486 9820
rect 15422 9760 15486 9764
rect 20610 9820 20674 9824
rect 20610 9764 20614 9820
rect 20614 9764 20670 9820
rect 20670 9764 20674 9820
rect 20610 9760 20674 9764
rect 20690 9820 20754 9824
rect 20690 9764 20694 9820
rect 20694 9764 20750 9820
rect 20750 9764 20754 9820
rect 20690 9760 20754 9764
rect 20770 9820 20834 9824
rect 20770 9764 20774 9820
rect 20774 9764 20830 9820
rect 20830 9764 20834 9820
rect 20770 9760 20834 9764
rect 20850 9820 20914 9824
rect 20850 9764 20854 9820
rect 20854 9764 20910 9820
rect 20910 9764 20914 9820
rect 20850 9760 20914 9764
rect 3666 9276 3730 9280
rect 3666 9220 3670 9276
rect 3670 9220 3726 9276
rect 3726 9220 3730 9276
rect 3666 9216 3730 9220
rect 3746 9276 3810 9280
rect 3746 9220 3750 9276
rect 3750 9220 3806 9276
rect 3806 9220 3810 9276
rect 3746 9216 3810 9220
rect 3826 9276 3890 9280
rect 3826 9220 3830 9276
rect 3830 9220 3886 9276
rect 3886 9220 3890 9276
rect 3826 9216 3890 9220
rect 3906 9276 3970 9280
rect 3906 9220 3910 9276
rect 3910 9220 3966 9276
rect 3966 9220 3970 9276
rect 3906 9216 3970 9220
rect 9094 9276 9158 9280
rect 9094 9220 9098 9276
rect 9098 9220 9154 9276
rect 9154 9220 9158 9276
rect 9094 9216 9158 9220
rect 9174 9276 9238 9280
rect 9174 9220 9178 9276
rect 9178 9220 9234 9276
rect 9234 9220 9238 9276
rect 9174 9216 9238 9220
rect 9254 9276 9318 9280
rect 9254 9220 9258 9276
rect 9258 9220 9314 9276
rect 9314 9220 9318 9276
rect 9254 9216 9318 9220
rect 9334 9276 9398 9280
rect 9334 9220 9338 9276
rect 9338 9220 9394 9276
rect 9394 9220 9398 9276
rect 9334 9216 9398 9220
rect 14522 9276 14586 9280
rect 14522 9220 14526 9276
rect 14526 9220 14582 9276
rect 14582 9220 14586 9276
rect 14522 9216 14586 9220
rect 14602 9276 14666 9280
rect 14602 9220 14606 9276
rect 14606 9220 14662 9276
rect 14662 9220 14666 9276
rect 14602 9216 14666 9220
rect 14682 9276 14746 9280
rect 14682 9220 14686 9276
rect 14686 9220 14742 9276
rect 14742 9220 14746 9276
rect 14682 9216 14746 9220
rect 14762 9276 14826 9280
rect 14762 9220 14766 9276
rect 14766 9220 14822 9276
rect 14822 9220 14826 9276
rect 14762 9216 14826 9220
rect 19950 9276 20014 9280
rect 19950 9220 19954 9276
rect 19954 9220 20010 9276
rect 20010 9220 20014 9276
rect 19950 9216 20014 9220
rect 20030 9276 20094 9280
rect 20030 9220 20034 9276
rect 20034 9220 20090 9276
rect 20090 9220 20094 9276
rect 20030 9216 20094 9220
rect 20110 9276 20174 9280
rect 20110 9220 20114 9276
rect 20114 9220 20170 9276
rect 20170 9220 20174 9276
rect 20110 9216 20174 9220
rect 20190 9276 20254 9280
rect 20190 9220 20194 9276
rect 20194 9220 20250 9276
rect 20250 9220 20254 9276
rect 20190 9216 20254 9220
rect 4326 8732 4390 8736
rect 4326 8676 4330 8732
rect 4330 8676 4386 8732
rect 4386 8676 4390 8732
rect 4326 8672 4390 8676
rect 4406 8732 4470 8736
rect 4406 8676 4410 8732
rect 4410 8676 4466 8732
rect 4466 8676 4470 8732
rect 4406 8672 4470 8676
rect 4486 8732 4550 8736
rect 4486 8676 4490 8732
rect 4490 8676 4546 8732
rect 4546 8676 4550 8732
rect 4486 8672 4550 8676
rect 4566 8732 4630 8736
rect 4566 8676 4570 8732
rect 4570 8676 4626 8732
rect 4626 8676 4630 8732
rect 4566 8672 4630 8676
rect 9754 8732 9818 8736
rect 9754 8676 9758 8732
rect 9758 8676 9814 8732
rect 9814 8676 9818 8732
rect 9754 8672 9818 8676
rect 9834 8732 9898 8736
rect 9834 8676 9838 8732
rect 9838 8676 9894 8732
rect 9894 8676 9898 8732
rect 9834 8672 9898 8676
rect 9914 8732 9978 8736
rect 9914 8676 9918 8732
rect 9918 8676 9974 8732
rect 9974 8676 9978 8732
rect 9914 8672 9978 8676
rect 9994 8732 10058 8736
rect 9994 8676 9998 8732
rect 9998 8676 10054 8732
rect 10054 8676 10058 8732
rect 9994 8672 10058 8676
rect 15182 8732 15246 8736
rect 15182 8676 15186 8732
rect 15186 8676 15242 8732
rect 15242 8676 15246 8732
rect 15182 8672 15246 8676
rect 15262 8732 15326 8736
rect 15262 8676 15266 8732
rect 15266 8676 15322 8732
rect 15322 8676 15326 8732
rect 15262 8672 15326 8676
rect 15342 8732 15406 8736
rect 15342 8676 15346 8732
rect 15346 8676 15402 8732
rect 15402 8676 15406 8732
rect 15342 8672 15406 8676
rect 15422 8732 15486 8736
rect 15422 8676 15426 8732
rect 15426 8676 15482 8732
rect 15482 8676 15486 8732
rect 15422 8672 15486 8676
rect 20610 8732 20674 8736
rect 20610 8676 20614 8732
rect 20614 8676 20670 8732
rect 20670 8676 20674 8732
rect 20610 8672 20674 8676
rect 20690 8732 20754 8736
rect 20690 8676 20694 8732
rect 20694 8676 20750 8732
rect 20750 8676 20754 8732
rect 20690 8672 20754 8676
rect 20770 8732 20834 8736
rect 20770 8676 20774 8732
rect 20774 8676 20830 8732
rect 20830 8676 20834 8732
rect 20770 8672 20834 8676
rect 20850 8732 20914 8736
rect 20850 8676 20854 8732
rect 20854 8676 20910 8732
rect 20910 8676 20914 8732
rect 20850 8672 20914 8676
rect 3666 8188 3730 8192
rect 3666 8132 3670 8188
rect 3670 8132 3726 8188
rect 3726 8132 3730 8188
rect 3666 8128 3730 8132
rect 3746 8188 3810 8192
rect 3746 8132 3750 8188
rect 3750 8132 3806 8188
rect 3806 8132 3810 8188
rect 3746 8128 3810 8132
rect 3826 8188 3890 8192
rect 3826 8132 3830 8188
rect 3830 8132 3886 8188
rect 3886 8132 3890 8188
rect 3826 8128 3890 8132
rect 3906 8188 3970 8192
rect 3906 8132 3910 8188
rect 3910 8132 3966 8188
rect 3966 8132 3970 8188
rect 3906 8128 3970 8132
rect 9094 8188 9158 8192
rect 9094 8132 9098 8188
rect 9098 8132 9154 8188
rect 9154 8132 9158 8188
rect 9094 8128 9158 8132
rect 9174 8188 9238 8192
rect 9174 8132 9178 8188
rect 9178 8132 9234 8188
rect 9234 8132 9238 8188
rect 9174 8128 9238 8132
rect 9254 8188 9318 8192
rect 9254 8132 9258 8188
rect 9258 8132 9314 8188
rect 9314 8132 9318 8188
rect 9254 8128 9318 8132
rect 9334 8188 9398 8192
rect 9334 8132 9338 8188
rect 9338 8132 9394 8188
rect 9394 8132 9398 8188
rect 9334 8128 9398 8132
rect 14522 8188 14586 8192
rect 14522 8132 14526 8188
rect 14526 8132 14582 8188
rect 14582 8132 14586 8188
rect 14522 8128 14586 8132
rect 14602 8188 14666 8192
rect 14602 8132 14606 8188
rect 14606 8132 14662 8188
rect 14662 8132 14666 8188
rect 14602 8128 14666 8132
rect 14682 8188 14746 8192
rect 14682 8132 14686 8188
rect 14686 8132 14742 8188
rect 14742 8132 14746 8188
rect 14682 8128 14746 8132
rect 14762 8188 14826 8192
rect 14762 8132 14766 8188
rect 14766 8132 14822 8188
rect 14822 8132 14826 8188
rect 14762 8128 14826 8132
rect 19950 8188 20014 8192
rect 19950 8132 19954 8188
rect 19954 8132 20010 8188
rect 20010 8132 20014 8188
rect 19950 8128 20014 8132
rect 20030 8188 20094 8192
rect 20030 8132 20034 8188
rect 20034 8132 20090 8188
rect 20090 8132 20094 8188
rect 20030 8128 20094 8132
rect 20110 8188 20174 8192
rect 20110 8132 20114 8188
rect 20114 8132 20170 8188
rect 20170 8132 20174 8188
rect 20110 8128 20174 8132
rect 20190 8188 20254 8192
rect 20190 8132 20194 8188
rect 20194 8132 20250 8188
rect 20250 8132 20254 8188
rect 20190 8128 20254 8132
rect 4326 7644 4390 7648
rect 4326 7588 4330 7644
rect 4330 7588 4386 7644
rect 4386 7588 4390 7644
rect 4326 7584 4390 7588
rect 4406 7644 4470 7648
rect 4406 7588 4410 7644
rect 4410 7588 4466 7644
rect 4466 7588 4470 7644
rect 4406 7584 4470 7588
rect 4486 7644 4550 7648
rect 4486 7588 4490 7644
rect 4490 7588 4546 7644
rect 4546 7588 4550 7644
rect 4486 7584 4550 7588
rect 4566 7644 4630 7648
rect 4566 7588 4570 7644
rect 4570 7588 4626 7644
rect 4626 7588 4630 7644
rect 4566 7584 4630 7588
rect 9754 7644 9818 7648
rect 9754 7588 9758 7644
rect 9758 7588 9814 7644
rect 9814 7588 9818 7644
rect 9754 7584 9818 7588
rect 9834 7644 9898 7648
rect 9834 7588 9838 7644
rect 9838 7588 9894 7644
rect 9894 7588 9898 7644
rect 9834 7584 9898 7588
rect 9914 7644 9978 7648
rect 9914 7588 9918 7644
rect 9918 7588 9974 7644
rect 9974 7588 9978 7644
rect 9914 7584 9978 7588
rect 9994 7644 10058 7648
rect 9994 7588 9998 7644
rect 9998 7588 10054 7644
rect 10054 7588 10058 7644
rect 9994 7584 10058 7588
rect 15182 7644 15246 7648
rect 15182 7588 15186 7644
rect 15186 7588 15242 7644
rect 15242 7588 15246 7644
rect 15182 7584 15246 7588
rect 15262 7644 15326 7648
rect 15262 7588 15266 7644
rect 15266 7588 15322 7644
rect 15322 7588 15326 7644
rect 15262 7584 15326 7588
rect 15342 7644 15406 7648
rect 15342 7588 15346 7644
rect 15346 7588 15402 7644
rect 15402 7588 15406 7644
rect 15342 7584 15406 7588
rect 15422 7644 15486 7648
rect 15422 7588 15426 7644
rect 15426 7588 15482 7644
rect 15482 7588 15486 7644
rect 15422 7584 15486 7588
rect 20610 7644 20674 7648
rect 20610 7588 20614 7644
rect 20614 7588 20670 7644
rect 20670 7588 20674 7644
rect 20610 7584 20674 7588
rect 20690 7644 20754 7648
rect 20690 7588 20694 7644
rect 20694 7588 20750 7644
rect 20750 7588 20754 7644
rect 20690 7584 20754 7588
rect 20770 7644 20834 7648
rect 20770 7588 20774 7644
rect 20774 7588 20830 7644
rect 20830 7588 20834 7644
rect 20770 7584 20834 7588
rect 20850 7644 20914 7648
rect 20850 7588 20854 7644
rect 20854 7588 20910 7644
rect 20910 7588 20914 7644
rect 20850 7584 20914 7588
rect 3666 7100 3730 7104
rect 3666 7044 3670 7100
rect 3670 7044 3726 7100
rect 3726 7044 3730 7100
rect 3666 7040 3730 7044
rect 3746 7100 3810 7104
rect 3746 7044 3750 7100
rect 3750 7044 3806 7100
rect 3806 7044 3810 7100
rect 3746 7040 3810 7044
rect 3826 7100 3890 7104
rect 3826 7044 3830 7100
rect 3830 7044 3886 7100
rect 3886 7044 3890 7100
rect 3826 7040 3890 7044
rect 3906 7100 3970 7104
rect 3906 7044 3910 7100
rect 3910 7044 3966 7100
rect 3966 7044 3970 7100
rect 3906 7040 3970 7044
rect 9094 7100 9158 7104
rect 9094 7044 9098 7100
rect 9098 7044 9154 7100
rect 9154 7044 9158 7100
rect 9094 7040 9158 7044
rect 9174 7100 9238 7104
rect 9174 7044 9178 7100
rect 9178 7044 9234 7100
rect 9234 7044 9238 7100
rect 9174 7040 9238 7044
rect 9254 7100 9318 7104
rect 9254 7044 9258 7100
rect 9258 7044 9314 7100
rect 9314 7044 9318 7100
rect 9254 7040 9318 7044
rect 9334 7100 9398 7104
rect 9334 7044 9338 7100
rect 9338 7044 9394 7100
rect 9394 7044 9398 7100
rect 9334 7040 9398 7044
rect 14522 7100 14586 7104
rect 14522 7044 14526 7100
rect 14526 7044 14582 7100
rect 14582 7044 14586 7100
rect 14522 7040 14586 7044
rect 14602 7100 14666 7104
rect 14602 7044 14606 7100
rect 14606 7044 14662 7100
rect 14662 7044 14666 7100
rect 14602 7040 14666 7044
rect 14682 7100 14746 7104
rect 14682 7044 14686 7100
rect 14686 7044 14742 7100
rect 14742 7044 14746 7100
rect 14682 7040 14746 7044
rect 14762 7100 14826 7104
rect 14762 7044 14766 7100
rect 14766 7044 14822 7100
rect 14822 7044 14826 7100
rect 14762 7040 14826 7044
rect 19950 7100 20014 7104
rect 19950 7044 19954 7100
rect 19954 7044 20010 7100
rect 20010 7044 20014 7100
rect 19950 7040 20014 7044
rect 20030 7100 20094 7104
rect 20030 7044 20034 7100
rect 20034 7044 20090 7100
rect 20090 7044 20094 7100
rect 20030 7040 20094 7044
rect 20110 7100 20174 7104
rect 20110 7044 20114 7100
rect 20114 7044 20170 7100
rect 20170 7044 20174 7100
rect 20110 7040 20174 7044
rect 20190 7100 20254 7104
rect 20190 7044 20194 7100
rect 20194 7044 20250 7100
rect 20250 7044 20254 7100
rect 20190 7040 20254 7044
rect 4326 6556 4390 6560
rect 4326 6500 4330 6556
rect 4330 6500 4386 6556
rect 4386 6500 4390 6556
rect 4326 6496 4390 6500
rect 4406 6556 4470 6560
rect 4406 6500 4410 6556
rect 4410 6500 4466 6556
rect 4466 6500 4470 6556
rect 4406 6496 4470 6500
rect 4486 6556 4550 6560
rect 4486 6500 4490 6556
rect 4490 6500 4546 6556
rect 4546 6500 4550 6556
rect 4486 6496 4550 6500
rect 4566 6556 4630 6560
rect 4566 6500 4570 6556
rect 4570 6500 4626 6556
rect 4626 6500 4630 6556
rect 4566 6496 4630 6500
rect 9754 6556 9818 6560
rect 9754 6500 9758 6556
rect 9758 6500 9814 6556
rect 9814 6500 9818 6556
rect 9754 6496 9818 6500
rect 9834 6556 9898 6560
rect 9834 6500 9838 6556
rect 9838 6500 9894 6556
rect 9894 6500 9898 6556
rect 9834 6496 9898 6500
rect 9914 6556 9978 6560
rect 9914 6500 9918 6556
rect 9918 6500 9974 6556
rect 9974 6500 9978 6556
rect 9914 6496 9978 6500
rect 9994 6556 10058 6560
rect 9994 6500 9998 6556
rect 9998 6500 10054 6556
rect 10054 6500 10058 6556
rect 9994 6496 10058 6500
rect 15182 6556 15246 6560
rect 15182 6500 15186 6556
rect 15186 6500 15242 6556
rect 15242 6500 15246 6556
rect 15182 6496 15246 6500
rect 15262 6556 15326 6560
rect 15262 6500 15266 6556
rect 15266 6500 15322 6556
rect 15322 6500 15326 6556
rect 15262 6496 15326 6500
rect 15342 6556 15406 6560
rect 15342 6500 15346 6556
rect 15346 6500 15402 6556
rect 15402 6500 15406 6556
rect 15342 6496 15406 6500
rect 15422 6556 15486 6560
rect 15422 6500 15426 6556
rect 15426 6500 15482 6556
rect 15482 6500 15486 6556
rect 15422 6496 15486 6500
rect 20610 6556 20674 6560
rect 20610 6500 20614 6556
rect 20614 6500 20670 6556
rect 20670 6500 20674 6556
rect 20610 6496 20674 6500
rect 20690 6556 20754 6560
rect 20690 6500 20694 6556
rect 20694 6500 20750 6556
rect 20750 6500 20754 6556
rect 20690 6496 20754 6500
rect 20770 6556 20834 6560
rect 20770 6500 20774 6556
rect 20774 6500 20830 6556
rect 20830 6500 20834 6556
rect 20770 6496 20834 6500
rect 20850 6556 20914 6560
rect 20850 6500 20854 6556
rect 20854 6500 20910 6556
rect 20910 6500 20914 6556
rect 20850 6496 20914 6500
rect 3666 6012 3730 6016
rect 3666 5956 3670 6012
rect 3670 5956 3726 6012
rect 3726 5956 3730 6012
rect 3666 5952 3730 5956
rect 3746 6012 3810 6016
rect 3746 5956 3750 6012
rect 3750 5956 3806 6012
rect 3806 5956 3810 6012
rect 3746 5952 3810 5956
rect 3826 6012 3890 6016
rect 3826 5956 3830 6012
rect 3830 5956 3886 6012
rect 3886 5956 3890 6012
rect 3826 5952 3890 5956
rect 3906 6012 3970 6016
rect 3906 5956 3910 6012
rect 3910 5956 3966 6012
rect 3966 5956 3970 6012
rect 3906 5952 3970 5956
rect 9094 6012 9158 6016
rect 9094 5956 9098 6012
rect 9098 5956 9154 6012
rect 9154 5956 9158 6012
rect 9094 5952 9158 5956
rect 9174 6012 9238 6016
rect 9174 5956 9178 6012
rect 9178 5956 9234 6012
rect 9234 5956 9238 6012
rect 9174 5952 9238 5956
rect 9254 6012 9318 6016
rect 9254 5956 9258 6012
rect 9258 5956 9314 6012
rect 9314 5956 9318 6012
rect 9254 5952 9318 5956
rect 9334 6012 9398 6016
rect 9334 5956 9338 6012
rect 9338 5956 9394 6012
rect 9394 5956 9398 6012
rect 9334 5952 9398 5956
rect 14522 6012 14586 6016
rect 14522 5956 14526 6012
rect 14526 5956 14582 6012
rect 14582 5956 14586 6012
rect 14522 5952 14586 5956
rect 14602 6012 14666 6016
rect 14602 5956 14606 6012
rect 14606 5956 14662 6012
rect 14662 5956 14666 6012
rect 14602 5952 14666 5956
rect 14682 6012 14746 6016
rect 14682 5956 14686 6012
rect 14686 5956 14742 6012
rect 14742 5956 14746 6012
rect 14682 5952 14746 5956
rect 14762 6012 14826 6016
rect 14762 5956 14766 6012
rect 14766 5956 14822 6012
rect 14822 5956 14826 6012
rect 14762 5952 14826 5956
rect 19950 6012 20014 6016
rect 19950 5956 19954 6012
rect 19954 5956 20010 6012
rect 20010 5956 20014 6012
rect 19950 5952 20014 5956
rect 20030 6012 20094 6016
rect 20030 5956 20034 6012
rect 20034 5956 20090 6012
rect 20090 5956 20094 6012
rect 20030 5952 20094 5956
rect 20110 6012 20174 6016
rect 20110 5956 20114 6012
rect 20114 5956 20170 6012
rect 20170 5956 20174 6012
rect 20110 5952 20174 5956
rect 20190 6012 20254 6016
rect 20190 5956 20194 6012
rect 20194 5956 20250 6012
rect 20250 5956 20254 6012
rect 20190 5952 20254 5956
rect 4326 5468 4390 5472
rect 4326 5412 4330 5468
rect 4330 5412 4386 5468
rect 4386 5412 4390 5468
rect 4326 5408 4390 5412
rect 4406 5468 4470 5472
rect 4406 5412 4410 5468
rect 4410 5412 4466 5468
rect 4466 5412 4470 5468
rect 4406 5408 4470 5412
rect 4486 5468 4550 5472
rect 4486 5412 4490 5468
rect 4490 5412 4546 5468
rect 4546 5412 4550 5468
rect 4486 5408 4550 5412
rect 4566 5468 4630 5472
rect 4566 5412 4570 5468
rect 4570 5412 4626 5468
rect 4626 5412 4630 5468
rect 4566 5408 4630 5412
rect 9754 5468 9818 5472
rect 9754 5412 9758 5468
rect 9758 5412 9814 5468
rect 9814 5412 9818 5468
rect 9754 5408 9818 5412
rect 9834 5468 9898 5472
rect 9834 5412 9838 5468
rect 9838 5412 9894 5468
rect 9894 5412 9898 5468
rect 9834 5408 9898 5412
rect 9914 5468 9978 5472
rect 9914 5412 9918 5468
rect 9918 5412 9974 5468
rect 9974 5412 9978 5468
rect 9914 5408 9978 5412
rect 9994 5468 10058 5472
rect 9994 5412 9998 5468
rect 9998 5412 10054 5468
rect 10054 5412 10058 5468
rect 9994 5408 10058 5412
rect 15182 5468 15246 5472
rect 15182 5412 15186 5468
rect 15186 5412 15242 5468
rect 15242 5412 15246 5468
rect 15182 5408 15246 5412
rect 15262 5468 15326 5472
rect 15262 5412 15266 5468
rect 15266 5412 15322 5468
rect 15322 5412 15326 5468
rect 15262 5408 15326 5412
rect 15342 5468 15406 5472
rect 15342 5412 15346 5468
rect 15346 5412 15402 5468
rect 15402 5412 15406 5468
rect 15342 5408 15406 5412
rect 15422 5468 15486 5472
rect 15422 5412 15426 5468
rect 15426 5412 15482 5468
rect 15482 5412 15486 5468
rect 15422 5408 15486 5412
rect 20610 5468 20674 5472
rect 20610 5412 20614 5468
rect 20614 5412 20670 5468
rect 20670 5412 20674 5468
rect 20610 5408 20674 5412
rect 20690 5468 20754 5472
rect 20690 5412 20694 5468
rect 20694 5412 20750 5468
rect 20750 5412 20754 5468
rect 20690 5408 20754 5412
rect 20770 5468 20834 5472
rect 20770 5412 20774 5468
rect 20774 5412 20830 5468
rect 20830 5412 20834 5468
rect 20770 5408 20834 5412
rect 20850 5468 20914 5472
rect 20850 5412 20854 5468
rect 20854 5412 20910 5468
rect 20910 5412 20914 5468
rect 20850 5408 20914 5412
rect 3666 4924 3730 4928
rect 3666 4868 3670 4924
rect 3670 4868 3726 4924
rect 3726 4868 3730 4924
rect 3666 4864 3730 4868
rect 3746 4924 3810 4928
rect 3746 4868 3750 4924
rect 3750 4868 3806 4924
rect 3806 4868 3810 4924
rect 3746 4864 3810 4868
rect 3826 4924 3890 4928
rect 3826 4868 3830 4924
rect 3830 4868 3886 4924
rect 3886 4868 3890 4924
rect 3826 4864 3890 4868
rect 3906 4924 3970 4928
rect 3906 4868 3910 4924
rect 3910 4868 3966 4924
rect 3966 4868 3970 4924
rect 3906 4864 3970 4868
rect 9094 4924 9158 4928
rect 9094 4868 9098 4924
rect 9098 4868 9154 4924
rect 9154 4868 9158 4924
rect 9094 4864 9158 4868
rect 9174 4924 9238 4928
rect 9174 4868 9178 4924
rect 9178 4868 9234 4924
rect 9234 4868 9238 4924
rect 9174 4864 9238 4868
rect 9254 4924 9318 4928
rect 9254 4868 9258 4924
rect 9258 4868 9314 4924
rect 9314 4868 9318 4924
rect 9254 4864 9318 4868
rect 9334 4924 9398 4928
rect 9334 4868 9338 4924
rect 9338 4868 9394 4924
rect 9394 4868 9398 4924
rect 9334 4864 9398 4868
rect 14522 4924 14586 4928
rect 14522 4868 14526 4924
rect 14526 4868 14582 4924
rect 14582 4868 14586 4924
rect 14522 4864 14586 4868
rect 14602 4924 14666 4928
rect 14602 4868 14606 4924
rect 14606 4868 14662 4924
rect 14662 4868 14666 4924
rect 14602 4864 14666 4868
rect 14682 4924 14746 4928
rect 14682 4868 14686 4924
rect 14686 4868 14742 4924
rect 14742 4868 14746 4924
rect 14682 4864 14746 4868
rect 14762 4924 14826 4928
rect 14762 4868 14766 4924
rect 14766 4868 14822 4924
rect 14822 4868 14826 4924
rect 14762 4864 14826 4868
rect 19950 4924 20014 4928
rect 19950 4868 19954 4924
rect 19954 4868 20010 4924
rect 20010 4868 20014 4924
rect 19950 4864 20014 4868
rect 20030 4924 20094 4928
rect 20030 4868 20034 4924
rect 20034 4868 20090 4924
rect 20090 4868 20094 4924
rect 20030 4864 20094 4868
rect 20110 4924 20174 4928
rect 20110 4868 20114 4924
rect 20114 4868 20170 4924
rect 20170 4868 20174 4924
rect 20110 4864 20174 4868
rect 20190 4924 20254 4928
rect 20190 4868 20194 4924
rect 20194 4868 20250 4924
rect 20250 4868 20254 4924
rect 20190 4864 20254 4868
rect 4326 4380 4390 4384
rect 4326 4324 4330 4380
rect 4330 4324 4386 4380
rect 4386 4324 4390 4380
rect 4326 4320 4390 4324
rect 4406 4380 4470 4384
rect 4406 4324 4410 4380
rect 4410 4324 4466 4380
rect 4466 4324 4470 4380
rect 4406 4320 4470 4324
rect 4486 4380 4550 4384
rect 4486 4324 4490 4380
rect 4490 4324 4546 4380
rect 4546 4324 4550 4380
rect 4486 4320 4550 4324
rect 4566 4380 4630 4384
rect 4566 4324 4570 4380
rect 4570 4324 4626 4380
rect 4626 4324 4630 4380
rect 4566 4320 4630 4324
rect 9754 4380 9818 4384
rect 9754 4324 9758 4380
rect 9758 4324 9814 4380
rect 9814 4324 9818 4380
rect 9754 4320 9818 4324
rect 9834 4380 9898 4384
rect 9834 4324 9838 4380
rect 9838 4324 9894 4380
rect 9894 4324 9898 4380
rect 9834 4320 9898 4324
rect 9914 4380 9978 4384
rect 9914 4324 9918 4380
rect 9918 4324 9974 4380
rect 9974 4324 9978 4380
rect 9914 4320 9978 4324
rect 9994 4380 10058 4384
rect 9994 4324 9998 4380
rect 9998 4324 10054 4380
rect 10054 4324 10058 4380
rect 9994 4320 10058 4324
rect 15182 4380 15246 4384
rect 15182 4324 15186 4380
rect 15186 4324 15242 4380
rect 15242 4324 15246 4380
rect 15182 4320 15246 4324
rect 15262 4380 15326 4384
rect 15262 4324 15266 4380
rect 15266 4324 15322 4380
rect 15322 4324 15326 4380
rect 15262 4320 15326 4324
rect 15342 4380 15406 4384
rect 15342 4324 15346 4380
rect 15346 4324 15402 4380
rect 15402 4324 15406 4380
rect 15342 4320 15406 4324
rect 15422 4380 15486 4384
rect 15422 4324 15426 4380
rect 15426 4324 15482 4380
rect 15482 4324 15486 4380
rect 15422 4320 15486 4324
rect 20610 4380 20674 4384
rect 20610 4324 20614 4380
rect 20614 4324 20670 4380
rect 20670 4324 20674 4380
rect 20610 4320 20674 4324
rect 20690 4380 20754 4384
rect 20690 4324 20694 4380
rect 20694 4324 20750 4380
rect 20750 4324 20754 4380
rect 20690 4320 20754 4324
rect 20770 4380 20834 4384
rect 20770 4324 20774 4380
rect 20774 4324 20830 4380
rect 20830 4324 20834 4380
rect 20770 4320 20834 4324
rect 20850 4380 20914 4384
rect 20850 4324 20854 4380
rect 20854 4324 20910 4380
rect 20910 4324 20914 4380
rect 20850 4320 20914 4324
rect 3666 3836 3730 3840
rect 3666 3780 3670 3836
rect 3670 3780 3726 3836
rect 3726 3780 3730 3836
rect 3666 3776 3730 3780
rect 3746 3836 3810 3840
rect 3746 3780 3750 3836
rect 3750 3780 3806 3836
rect 3806 3780 3810 3836
rect 3746 3776 3810 3780
rect 3826 3836 3890 3840
rect 3826 3780 3830 3836
rect 3830 3780 3886 3836
rect 3886 3780 3890 3836
rect 3826 3776 3890 3780
rect 3906 3836 3970 3840
rect 3906 3780 3910 3836
rect 3910 3780 3966 3836
rect 3966 3780 3970 3836
rect 3906 3776 3970 3780
rect 9094 3836 9158 3840
rect 9094 3780 9098 3836
rect 9098 3780 9154 3836
rect 9154 3780 9158 3836
rect 9094 3776 9158 3780
rect 9174 3836 9238 3840
rect 9174 3780 9178 3836
rect 9178 3780 9234 3836
rect 9234 3780 9238 3836
rect 9174 3776 9238 3780
rect 9254 3836 9318 3840
rect 9254 3780 9258 3836
rect 9258 3780 9314 3836
rect 9314 3780 9318 3836
rect 9254 3776 9318 3780
rect 9334 3836 9398 3840
rect 9334 3780 9338 3836
rect 9338 3780 9394 3836
rect 9394 3780 9398 3836
rect 9334 3776 9398 3780
rect 14522 3836 14586 3840
rect 14522 3780 14526 3836
rect 14526 3780 14582 3836
rect 14582 3780 14586 3836
rect 14522 3776 14586 3780
rect 14602 3836 14666 3840
rect 14602 3780 14606 3836
rect 14606 3780 14662 3836
rect 14662 3780 14666 3836
rect 14602 3776 14666 3780
rect 14682 3836 14746 3840
rect 14682 3780 14686 3836
rect 14686 3780 14742 3836
rect 14742 3780 14746 3836
rect 14682 3776 14746 3780
rect 14762 3836 14826 3840
rect 14762 3780 14766 3836
rect 14766 3780 14822 3836
rect 14822 3780 14826 3836
rect 14762 3776 14826 3780
rect 19950 3836 20014 3840
rect 19950 3780 19954 3836
rect 19954 3780 20010 3836
rect 20010 3780 20014 3836
rect 19950 3776 20014 3780
rect 20030 3836 20094 3840
rect 20030 3780 20034 3836
rect 20034 3780 20090 3836
rect 20090 3780 20094 3836
rect 20030 3776 20094 3780
rect 20110 3836 20174 3840
rect 20110 3780 20114 3836
rect 20114 3780 20170 3836
rect 20170 3780 20174 3836
rect 20110 3776 20174 3780
rect 20190 3836 20254 3840
rect 20190 3780 20194 3836
rect 20194 3780 20250 3836
rect 20250 3780 20254 3836
rect 20190 3776 20254 3780
rect 4326 3292 4390 3296
rect 4326 3236 4330 3292
rect 4330 3236 4386 3292
rect 4386 3236 4390 3292
rect 4326 3232 4390 3236
rect 4406 3292 4470 3296
rect 4406 3236 4410 3292
rect 4410 3236 4466 3292
rect 4466 3236 4470 3292
rect 4406 3232 4470 3236
rect 4486 3292 4550 3296
rect 4486 3236 4490 3292
rect 4490 3236 4546 3292
rect 4546 3236 4550 3292
rect 4486 3232 4550 3236
rect 4566 3292 4630 3296
rect 4566 3236 4570 3292
rect 4570 3236 4626 3292
rect 4626 3236 4630 3292
rect 4566 3232 4630 3236
rect 9754 3292 9818 3296
rect 9754 3236 9758 3292
rect 9758 3236 9814 3292
rect 9814 3236 9818 3292
rect 9754 3232 9818 3236
rect 9834 3292 9898 3296
rect 9834 3236 9838 3292
rect 9838 3236 9894 3292
rect 9894 3236 9898 3292
rect 9834 3232 9898 3236
rect 9914 3292 9978 3296
rect 9914 3236 9918 3292
rect 9918 3236 9974 3292
rect 9974 3236 9978 3292
rect 9914 3232 9978 3236
rect 9994 3292 10058 3296
rect 9994 3236 9998 3292
rect 9998 3236 10054 3292
rect 10054 3236 10058 3292
rect 9994 3232 10058 3236
rect 15182 3292 15246 3296
rect 15182 3236 15186 3292
rect 15186 3236 15242 3292
rect 15242 3236 15246 3292
rect 15182 3232 15246 3236
rect 15262 3292 15326 3296
rect 15262 3236 15266 3292
rect 15266 3236 15322 3292
rect 15322 3236 15326 3292
rect 15262 3232 15326 3236
rect 15342 3292 15406 3296
rect 15342 3236 15346 3292
rect 15346 3236 15402 3292
rect 15402 3236 15406 3292
rect 15342 3232 15406 3236
rect 15422 3292 15486 3296
rect 15422 3236 15426 3292
rect 15426 3236 15482 3292
rect 15482 3236 15486 3292
rect 15422 3232 15486 3236
rect 20610 3292 20674 3296
rect 20610 3236 20614 3292
rect 20614 3236 20670 3292
rect 20670 3236 20674 3292
rect 20610 3232 20674 3236
rect 20690 3292 20754 3296
rect 20690 3236 20694 3292
rect 20694 3236 20750 3292
rect 20750 3236 20754 3292
rect 20690 3232 20754 3236
rect 20770 3292 20834 3296
rect 20770 3236 20774 3292
rect 20774 3236 20830 3292
rect 20830 3236 20834 3292
rect 20770 3232 20834 3236
rect 20850 3292 20914 3296
rect 20850 3236 20854 3292
rect 20854 3236 20910 3292
rect 20910 3236 20914 3292
rect 20850 3232 20914 3236
rect 3666 2748 3730 2752
rect 3666 2692 3670 2748
rect 3670 2692 3726 2748
rect 3726 2692 3730 2748
rect 3666 2688 3730 2692
rect 3746 2748 3810 2752
rect 3746 2692 3750 2748
rect 3750 2692 3806 2748
rect 3806 2692 3810 2748
rect 3746 2688 3810 2692
rect 3826 2748 3890 2752
rect 3826 2692 3830 2748
rect 3830 2692 3886 2748
rect 3886 2692 3890 2748
rect 3826 2688 3890 2692
rect 3906 2748 3970 2752
rect 3906 2692 3910 2748
rect 3910 2692 3966 2748
rect 3966 2692 3970 2748
rect 3906 2688 3970 2692
rect 9094 2748 9158 2752
rect 9094 2692 9098 2748
rect 9098 2692 9154 2748
rect 9154 2692 9158 2748
rect 9094 2688 9158 2692
rect 9174 2748 9238 2752
rect 9174 2692 9178 2748
rect 9178 2692 9234 2748
rect 9234 2692 9238 2748
rect 9174 2688 9238 2692
rect 9254 2748 9318 2752
rect 9254 2692 9258 2748
rect 9258 2692 9314 2748
rect 9314 2692 9318 2748
rect 9254 2688 9318 2692
rect 9334 2748 9398 2752
rect 9334 2692 9338 2748
rect 9338 2692 9394 2748
rect 9394 2692 9398 2748
rect 9334 2688 9398 2692
rect 14522 2748 14586 2752
rect 14522 2692 14526 2748
rect 14526 2692 14582 2748
rect 14582 2692 14586 2748
rect 14522 2688 14586 2692
rect 14602 2748 14666 2752
rect 14602 2692 14606 2748
rect 14606 2692 14662 2748
rect 14662 2692 14666 2748
rect 14602 2688 14666 2692
rect 14682 2748 14746 2752
rect 14682 2692 14686 2748
rect 14686 2692 14742 2748
rect 14742 2692 14746 2748
rect 14682 2688 14746 2692
rect 14762 2748 14826 2752
rect 14762 2692 14766 2748
rect 14766 2692 14822 2748
rect 14822 2692 14826 2748
rect 14762 2688 14826 2692
rect 19950 2748 20014 2752
rect 19950 2692 19954 2748
rect 19954 2692 20010 2748
rect 20010 2692 20014 2748
rect 19950 2688 20014 2692
rect 20030 2748 20094 2752
rect 20030 2692 20034 2748
rect 20034 2692 20090 2748
rect 20090 2692 20094 2748
rect 20030 2688 20094 2692
rect 20110 2748 20174 2752
rect 20110 2692 20114 2748
rect 20114 2692 20170 2748
rect 20170 2692 20174 2748
rect 20110 2688 20174 2692
rect 20190 2748 20254 2752
rect 20190 2692 20194 2748
rect 20194 2692 20250 2748
rect 20250 2692 20254 2748
rect 20190 2688 20254 2692
rect 4326 2204 4390 2208
rect 4326 2148 4330 2204
rect 4330 2148 4386 2204
rect 4386 2148 4390 2204
rect 4326 2144 4390 2148
rect 4406 2204 4470 2208
rect 4406 2148 4410 2204
rect 4410 2148 4466 2204
rect 4466 2148 4470 2204
rect 4406 2144 4470 2148
rect 4486 2204 4550 2208
rect 4486 2148 4490 2204
rect 4490 2148 4546 2204
rect 4546 2148 4550 2204
rect 4486 2144 4550 2148
rect 4566 2204 4630 2208
rect 4566 2148 4570 2204
rect 4570 2148 4626 2204
rect 4626 2148 4630 2204
rect 4566 2144 4630 2148
rect 9754 2204 9818 2208
rect 9754 2148 9758 2204
rect 9758 2148 9814 2204
rect 9814 2148 9818 2204
rect 9754 2144 9818 2148
rect 9834 2204 9898 2208
rect 9834 2148 9838 2204
rect 9838 2148 9894 2204
rect 9894 2148 9898 2204
rect 9834 2144 9898 2148
rect 9914 2204 9978 2208
rect 9914 2148 9918 2204
rect 9918 2148 9974 2204
rect 9974 2148 9978 2204
rect 9914 2144 9978 2148
rect 9994 2204 10058 2208
rect 9994 2148 9998 2204
rect 9998 2148 10054 2204
rect 10054 2148 10058 2204
rect 9994 2144 10058 2148
rect 15182 2204 15246 2208
rect 15182 2148 15186 2204
rect 15186 2148 15242 2204
rect 15242 2148 15246 2204
rect 15182 2144 15246 2148
rect 15262 2204 15326 2208
rect 15262 2148 15266 2204
rect 15266 2148 15322 2204
rect 15322 2148 15326 2204
rect 15262 2144 15326 2148
rect 15342 2204 15406 2208
rect 15342 2148 15346 2204
rect 15346 2148 15402 2204
rect 15402 2148 15406 2204
rect 15342 2144 15406 2148
rect 15422 2204 15486 2208
rect 15422 2148 15426 2204
rect 15426 2148 15482 2204
rect 15482 2148 15486 2204
rect 15422 2144 15486 2148
rect 20610 2204 20674 2208
rect 20610 2148 20614 2204
rect 20614 2148 20670 2204
rect 20670 2148 20674 2204
rect 20610 2144 20674 2148
rect 20690 2204 20754 2208
rect 20690 2148 20694 2204
rect 20694 2148 20750 2204
rect 20750 2148 20754 2204
rect 20690 2144 20754 2148
rect 20770 2204 20834 2208
rect 20770 2148 20774 2204
rect 20774 2148 20830 2204
rect 20830 2148 20834 2204
rect 20770 2144 20834 2148
rect 20850 2204 20914 2208
rect 20850 2148 20854 2204
rect 20854 2148 20910 2204
rect 20910 2148 20914 2204
rect 20850 2144 20914 2148
<< metal4 >>
rect 3658 21248 3978 21808
rect 3658 21184 3666 21248
rect 3730 21184 3746 21248
rect 3810 21184 3826 21248
rect 3890 21184 3906 21248
rect 3970 21184 3978 21248
rect 3658 20160 3978 21184
rect 3658 20096 3666 20160
rect 3730 20096 3746 20160
rect 3810 20096 3826 20160
rect 3890 20096 3906 20160
rect 3970 20096 3978 20160
rect 3658 19430 3978 20096
rect 3658 19194 3700 19430
rect 3936 19194 3978 19430
rect 3658 19072 3978 19194
rect 3658 19008 3666 19072
rect 3730 19008 3746 19072
rect 3810 19008 3826 19072
rect 3890 19008 3906 19072
rect 3970 19008 3978 19072
rect 3658 17984 3978 19008
rect 3658 17920 3666 17984
rect 3730 17920 3746 17984
rect 3810 17920 3826 17984
rect 3890 17920 3906 17984
rect 3970 17920 3978 17984
rect 3658 16896 3978 17920
rect 3658 16832 3666 16896
rect 3730 16832 3746 16896
rect 3810 16832 3826 16896
rect 3890 16832 3906 16896
rect 3970 16832 3978 16896
rect 3658 15808 3978 16832
rect 3658 15744 3666 15808
rect 3730 15744 3746 15808
rect 3810 15744 3826 15808
rect 3890 15744 3906 15808
rect 3970 15744 3978 15808
rect 3658 14720 3978 15744
rect 3658 14656 3666 14720
rect 3730 14656 3746 14720
rect 3810 14656 3826 14720
rect 3890 14656 3906 14720
rect 3970 14656 3978 14720
rect 3658 14534 3978 14656
rect 3658 14298 3700 14534
rect 3936 14298 3978 14534
rect 3658 13632 3978 14298
rect 3658 13568 3666 13632
rect 3730 13568 3746 13632
rect 3810 13568 3826 13632
rect 3890 13568 3906 13632
rect 3970 13568 3978 13632
rect 3658 12544 3978 13568
rect 3658 12480 3666 12544
rect 3730 12480 3746 12544
rect 3810 12480 3826 12544
rect 3890 12480 3906 12544
rect 3970 12480 3978 12544
rect 3658 11456 3978 12480
rect 3658 11392 3666 11456
rect 3730 11392 3746 11456
rect 3810 11392 3826 11456
rect 3890 11392 3906 11456
rect 3970 11392 3978 11456
rect 3658 10368 3978 11392
rect 3658 10304 3666 10368
rect 3730 10304 3746 10368
rect 3810 10304 3826 10368
rect 3890 10304 3906 10368
rect 3970 10304 3978 10368
rect 3658 9638 3978 10304
rect 3658 9402 3700 9638
rect 3936 9402 3978 9638
rect 3658 9280 3978 9402
rect 3658 9216 3666 9280
rect 3730 9216 3746 9280
rect 3810 9216 3826 9280
rect 3890 9216 3906 9280
rect 3970 9216 3978 9280
rect 3658 8192 3978 9216
rect 3658 8128 3666 8192
rect 3730 8128 3746 8192
rect 3810 8128 3826 8192
rect 3890 8128 3906 8192
rect 3970 8128 3978 8192
rect 3658 7104 3978 8128
rect 3658 7040 3666 7104
rect 3730 7040 3746 7104
rect 3810 7040 3826 7104
rect 3890 7040 3906 7104
rect 3970 7040 3978 7104
rect 3658 6016 3978 7040
rect 3658 5952 3666 6016
rect 3730 5952 3746 6016
rect 3810 5952 3826 6016
rect 3890 5952 3906 6016
rect 3970 5952 3978 6016
rect 3658 4928 3978 5952
rect 3658 4864 3666 4928
rect 3730 4864 3746 4928
rect 3810 4864 3826 4928
rect 3890 4864 3906 4928
rect 3970 4864 3978 4928
rect 3658 4742 3978 4864
rect 3658 4506 3700 4742
rect 3936 4506 3978 4742
rect 3658 3840 3978 4506
rect 3658 3776 3666 3840
rect 3730 3776 3746 3840
rect 3810 3776 3826 3840
rect 3890 3776 3906 3840
rect 3970 3776 3978 3840
rect 3658 2752 3978 3776
rect 3658 2688 3666 2752
rect 3730 2688 3746 2752
rect 3810 2688 3826 2752
rect 3890 2688 3906 2752
rect 3970 2688 3978 2752
rect 3658 2128 3978 2688
rect 4318 21792 4638 21808
rect 4318 21728 4326 21792
rect 4390 21728 4406 21792
rect 4470 21728 4486 21792
rect 4550 21728 4566 21792
rect 4630 21728 4638 21792
rect 4318 20704 4638 21728
rect 4318 20640 4326 20704
rect 4390 20640 4406 20704
rect 4470 20640 4486 20704
rect 4550 20640 4566 20704
rect 4630 20640 4638 20704
rect 4318 20090 4638 20640
rect 4318 19854 4360 20090
rect 4596 19854 4638 20090
rect 4318 19616 4638 19854
rect 4318 19552 4326 19616
rect 4390 19552 4406 19616
rect 4470 19552 4486 19616
rect 4550 19552 4566 19616
rect 4630 19552 4638 19616
rect 4318 18528 4638 19552
rect 4318 18464 4326 18528
rect 4390 18464 4406 18528
rect 4470 18464 4486 18528
rect 4550 18464 4566 18528
rect 4630 18464 4638 18528
rect 4318 17440 4638 18464
rect 4318 17376 4326 17440
rect 4390 17376 4406 17440
rect 4470 17376 4486 17440
rect 4550 17376 4566 17440
rect 4630 17376 4638 17440
rect 4318 16352 4638 17376
rect 4318 16288 4326 16352
rect 4390 16288 4406 16352
rect 4470 16288 4486 16352
rect 4550 16288 4566 16352
rect 4630 16288 4638 16352
rect 4318 15264 4638 16288
rect 4318 15200 4326 15264
rect 4390 15200 4406 15264
rect 4470 15200 4486 15264
rect 4550 15200 4566 15264
rect 4630 15200 4638 15264
rect 4318 15194 4638 15200
rect 4318 14958 4360 15194
rect 4596 14958 4638 15194
rect 4318 14176 4638 14958
rect 4318 14112 4326 14176
rect 4390 14112 4406 14176
rect 4470 14112 4486 14176
rect 4550 14112 4566 14176
rect 4630 14112 4638 14176
rect 4318 13088 4638 14112
rect 4318 13024 4326 13088
rect 4390 13024 4406 13088
rect 4470 13024 4486 13088
rect 4550 13024 4566 13088
rect 4630 13024 4638 13088
rect 4318 12000 4638 13024
rect 4318 11936 4326 12000
rect 4390 11936 4406 12000
rect 4470 11936 4486 12000
rect 4550 11936 4566 12000
rect 4630 11936 4638 12000
rect 4318 10912 4638 11936
rect 4318 10848 4326 10912
rect 4390 10848 4406 10912
rect 4470 10848 4486 10912
rect 4550 10848 4566 10912
rect 4630 10848 4638 10912
rect 4318 10298 4638 10848
rect 4318 10062 4360 10298
rect 4596 10062 4638 10298
rect 4318 9824 4638 10062
rect 4318 9760 4326 9824
rect 4390 9760 4406 9824
rect 4470 9760 4486 9824
rect 4550 9760 4566 9824
rect 4630 9760 4638 9824
rect 4318 8736 4638 9760
rect 4318 8672 4326 8736
rect 4390 8672 4406 8736
rect 4470 8672 4486 8736
rect 4550 8672 4566 8736
rect 4630 8672 4638 8736
rect 4318 7648 4638 8672
rect 4318 7584 4326 7648
rect 4390 7584 4406 7648
rect 4470 7584 4486 7648
rect 4550 7584 4566 7648
rect 4630 7584 4638 7648
rect 4318 6560 4638 7584
rect 4318 6496 4326 6560
rect 4390 6496 4406 6560
rect 4470 6496 4486 6560
rect 4550 6496 4566 6560
rect 4630 6496 4638 6560
rect 4318 5472 4638 6496
rect 4318 5408 4326 5472
rect 4390 5408 4406 5472
rect 4470 5408 4486 5472
rect 4550 5408 4566 5472
rect 4630 5408 4638 5472
rect 4318 5402 4638 5408
rect 4318 5166 4360 5402
rect 4596 5166 4638 5402
rect 4318 4384 4638 5166
rect 4318 4320 4326 4384
rect 4390 4320 4406 4384
rect 4470 4320 4486 4384
rect 4550 4320 4566 4384
rect 4630 4320 4638 4384
rect 4318 3296 4638 4320
rect 4318 3232 4326 3296
rect 4390 3232 4406 3296
rect 4470 3232 4486 3296
rect 4550 3232 4566 3296
rect 4630 3232 4638 3296
rect 4318 2208 4638 3232
rect 4318 2144 4326 2208
rect 4390 2144 4406 2208
rect 4470 2144 4486 2208
rect 4550 2144 4566 2208
rect 4630 2144 4638 2208
rect 4318 2128 4638 2144
rect 9086 21248 9406 21808
rect 9086 21184 9094 21248
rect 9158 21184 9174 21248
rect 9238 21184 9254 21248
rect 9318 21184 9334 21248
rect 9398 21184 9406 21248
rect 9086 20160 9406 21184
rect 9086 20096 9094 20160
rect 9158 20096 9174 20160
rect 9238 20096 9254 20160
rect 9318 20096 9334 20160
rect 9398 20096 9406 20160
rect 9086 19430 9406 20096
rect 9086 19194 9128 19430
rect 9364 19194 9406 19430
rect 9086 19072 9406 19194
rect 9086 19008 9094 19072
rect 9158 19008 9174 19072
rect 9238 19008 9254 19072
rect 9318 19008 9334 19072
rect 9398 19008 9406 19072
rect 9086 17984 9406 19008
rect 9086 17920 9094 17984
rect 9158 17920 9174 17984
rect 9238 17920 9254 17984
rect 9318 17920 9334 17984
rect 9398 17920 9406 17984
rect 9086 16896 9406 17920
rect 9086 16832 9094 16896
rect 9158 16832 9174 16896
rect 9238 16832 9254 16896
rect 9318 16832 9334 16896
rect 9398 16832 9406 16896
rect 9086 15808 9406 16832
rect 9086 15744 9094 15808
rect 9158 15744 9174 15808
rect 9238 15744 9254 15808
rect 9318 15744 9334 15808
rect 9398 15744 9406 15808
rect 9086 14720 9406 15744
rect 9086 14656 9094 14720
rect 9158 14656 9174 14720
rect 9238 14656 9254 14720
rect 9318 14656 9334 14720
rect 9398 14656 9406 14720
rect 9086 14534 9406 14656
rect 9086 14298 9128 14534
rect 9364 14298 9406 14534
rect 9086 13632 9406 14298
rect 9086 13568 9094 13632
rect 9158 13568 9174 13632
rect 9238 13568 9254 13632
rect 9318 13568 9334 13632
rect 9398 13568 9406 13632
rect 9086 12544 9406 13568
rect 9086 12480 9094 12544
rect 9158 12480 9174 12544
rect 9238 12480 9254 12544
rect 9318 12480 9334 12544
rect 9398 12480 9406 12544
rect 9086 11456 9406 12480
rect 9086 11392 9094 11456
rect 9158 11392 9174 11456
rect 9238 11392 9254 11456
rect 9318 11392 9334 11456
rect 9398 11392 9406 11456
rect 9086 10368 9406 11392
rect 9086 10304 9094 10368
rect 9158 10304 9174 10368
rect 9238 10304 9254 10368
rect 9318 10304 9334 10368
rect 9398 10304 9406 10368
rect 9086 9638 9406 10304
rect 9086 9402 9128 9638
rect 9364 9402 9406 9638
rect 9086 9280 9406 9402
rect 9086 9216 9094 9280
rect 9158 9216 9174 9280
rect 9238 9216 9254 9280
rect 9318 9216 9334 9280
rect 9398 9216 9406 9280
rect 9086 8192 9406 9216
rect 9086 8128 9094 8192
rect 9158 8128 9174 8192
rect 9238 8128 9254 8192
rect 9318 8128 9334 8192
rect 9398 8128 9406 8192
rect 9086 7104 9406 8128
rect 9086 7040 9094 7104
rect 9158 7040 9174 7104
rect 9238 7040 9254 7104
rect 9318 7040 9334 7104
rect 9398 7040 9406 7104
rect 9086 6016 9406 7040
rect 9086 5952 9094 6016
rect 9158 5952 9174 6016
rect 9238 5952 9254 6016
rect 9318 5952 9334 6016
rect 9398 5952 9406 6016
rect 9086 4928 9406 5952
rect 9086 4864 9094 4928
rect 9158 4864 9174 4928
rect 9238 4864 9254 4928
rect 9318 4864 9334 4928
rect 9398 4864 9406 4928
rect 9086 4742 9406 4864
rect 9086 4506 9128 4742
rect 9364 4506 9406 4742
rect 9086 3840 9406 4506
rect 9086 3776 9094 3840
rect 9158 3776 9174 3840
rect 9238 3776 9254 3840
rect 9318 3776 9334 3840
rect 9398 3776 9406 3840
rect 9086 2752 9406 3776
rect 9086 2688 9094 2752
rect 9158 2688 9174 2752
rect 9238 2688 9254 2752
rect 9318 2688 9334 2752
rect 9398 2688 9406 2752
rect 9086 2128 9406 2688
rect 9746 21792 10066 21808
rect 9746 21728 9754 21792
rect 9818 21728 9834 21792
rect 9898 21728 9914 21792
rect 9978 21728 9994 21792
rect 10058 21728 10066 21792
rect 9746 20704 10066 21728
rect 9746 20640 9754 20704
rect 9818 20640 9834 20704
rect 9898 20640 9914 20704
rect 9978 20640 9994 20704
rect 10058 20640 10066 20704
rect 9746 20090 10066 20640
rect 9746 19854 9788 20090
rect 10024 19854 10066 20090
rect 9746 19616 10066 19854
rect 9746 19552 9754 19616
rect 9818 19552 9834 19616
rect 9898 19552 9914 19616
rect 9978 19552 9994 19616
rect 10058 19552 10066 19616
rect 9746 18528 10066 19552
rect 9746 18464 9754 18528
rect 9818 18464 9834 18528
rect 9898 18464 9914 18528
rect 9978 18464 9994 18528
rect 10058 18464 10066 18528
rect 9746 17440 10066 18464
rect 9746 17376 9754 17440
rect 9818 17376 9834 17440
rect 9898 17376 9914 17440
rect 9978 17376 9994 17440
rect 10058 17376 10066 17440
rect 9746 16352 10066 17376
rect 9746 16288 9754 16352
rect 9818 16288 9834 16352
rect 9898 16288 9914 16352
rect 9978 16288 9994 16352
rect 10058 16288 10066 16352
rect 9746 15264 10066 16288
rect 9746 15200 9754 15264
rect 9818 15200 9834 15264
rect 9898 15200 9914 15264
rect 9978 15200 9994 15264
rect 10058 15200 10066 15264
rect 9746 15194 10066 15200
rect 9746 14958 9788 15194
rect 10024 14958 10066 15194
rect 9746 14176 10066 14958
rect 9746 14112 9754 14176
rect 9818 14112 9834 14176
rect 9898 14112 9914 14176
rect 9978 14112 9994 14176
rect 10058 14112 10066 14176
rect 9746 13088 10066 14112
rect 9746 13024 9754 13088
rect 9818 13024 9834 13088
rect 9898 13024 9914 13088
rect 9978 13024 9994 13088
rect 10058 13024 10066 13088
rect 9746 12000 10066 13024
rect 9746 11936 9754 12000
rect 9818 11936 9834 12000
rect 9898 11936 9914 12000
rect 9978 11936 9994 12000
rect 10058 11936 10066 12000
rect 9746 10912 10066 11936
rect 9746 10848 9754 10912
rect 9818 10848 9834 10912
rect 9898 10848 9914 10912
rect 9978 10848 9994 10912
rect 10058 10848 10066 10912
rect 9746 10298 10066 10848
rect 9746 10062 9788 10298
rect 10024 10062 10066 10298
rect 9746 9824 10066 10062
rect 9746 9760 9754 9824
rect 9818 9760 9834 9824
rect 9898 9760 9914 9824
rect 9978 9760 9994 9824
rect 10058 9760 10066 9824
rect 9746 8736 10066 9760
rect 9746 8672 9754 8736
rect 9818 8672 9834 8736
rect 9898 8672 9914 8736
rect 9978 8672 9994 8736
rect 10058 8672 10066 8736
rect 9746 7648 10066 8672
rect 9746 7584 9754 7648
rect 9818 7584 9834 7648
rect 9898 7584 9914 7648
rect 9978 7584 9994 7648
rect 10058 7584 10066 7648
rect 9746 6560 10066 7584
rect 9746 6496 9754 6560
rect 9818 6496 9834 6560
rect 9898 6496 9914 6560
rect 9978 6496 9994 6560
rect 10058 6496 10066 6560
rect 9746 5472 10066 6496
rect 9746 5408 9754 5472
rect 9818 5408 9834 5472
rect 9898 5408 9914 5472
rect 9978 5408 9994 5472
rect 10058 5408 10066 5472
rect 9746 5402 10066 5408
rect 9746 5166 9788 5402
rect 10024 5166 10066 5402
rect 9746 4384 10066 5166
rect 9746 4320 9754 4384
rect 9818 4320 9834 4384
rect 9898 4320 9914 4384
rect 9978 4320 9994 4384
rect 10058 4320 10066 4384
rect 9746 3296 10066 4320
rect 9746 3232 9754 3296
rect 9818 3232 9834 3296
rect 9898 3232 9914 3296
rect 9978 3232 9994 3296
rect 10058 3232 10066 3296
rect 9746 2208 10066 3232
rect 9746 2144 9754 2208
rect 9818 2144 9834 2208
rect 9898 2144 9914 2208
rect 9978 2144 9994 2208
rect 10058 2144 10066 2208
rect 9746 2128 10066 2144
rect 14514 21248 14834 21808
rect 14514 21184 14522 21248
rect 14586 21184 14602 21248
rect 14666 21184 14682 21248
rect 14746 21184 14762 21248
rect 14826 21184 14834 21248
rect 14514 20160 14834 21184
rect 14514 20096 14522 20160
rect 14586 20096 14602 20160
rect 14666 20096 14682 20160
rect 14746 20096 14762 20160
rect 14826 20096 14834 20160
rect 14514 19430 14834 20096
rect 14514 19194 14556 19430
rect 14792 19194 14834 19430
rect 14514 19072 14834 19194
rect 14514 19008 14522 19072
rect 14586 19008 14602 19072
rect 14666 19008 14682 19072
rect 14746 19008 14762 19072
rect 14826 19008 14834 19072
rect 14514 17984 14834 19008
rect 14514 17920 14522 17984
rect 14586 17920 14602 17984
rect 14666 17920 14682 17984
rect 14746 17920 14762 17984
rect 14826 17920 14834 17984
rect 14514 16896 14834 17920
rect 14514 16832 14522 16896
rect 14586 16832 14602 16896
rect 14666 16832 14682 16896
rect 14746 16832 14762 16896
rect 14826 16832 14834 16896
rect 14514 15808 14834 16832
rect 14514 15744 14522 15808
rect 14586 15744 14602 15808
rect 14666 15744 14682 15808
rect 14746 15744 14762 15808
rect 14826 15744 14834 15808
rect 14514 14720 14834 15744
rect 14514 14656 14522 14720
rect 14586 14656 14602 14720
rect 14666 14656 14682 14720
rect 14746 14656 14762 14720
rect 14826 14656 14834 14720
rect 14514 14534 14834 14656
rect 14514 14298 14556 14534
rect 14792 14298 14834 14534
rect 14514 13632 14834 14298
rect 14514 13568 14522 13632
rect 14586 13568 14602 13632
rect 14666 13568 14682 13632
rect 14746 13568 14762 13632
rect 14826 13568 14834 13632
rect 14514 12544 14834 13568
rect 14514 12480 14522 12544
rect 14586 12480 14602 12544
rect 14666 12480 14682 12544
rect 14746 12480 14762 12544
rect 14826 12480 14834 12544
rect 14514 11456 14834 12480
rect 14514 11392 14522 11456
rect 14586 11392 14602 11456
rect 14666 11392 14682 11456
rect 14746 11392 14762 11456
rect 14826 11392 14834 11456
rect 14514 10368 14834 11392
rect 14514 10304 14522 10368
rect 14586 10304 14602 10368
rect 14666 10304 14682 10368
rect 14746 10304 14762 10368
rect 14826 10304 14834 10368
rect 14514 9638 14834 10304
rect 14514 9402 14556 9638
rect 14792 9402 14834 9638
rect 14514 9280 14834 9402
rect 14514 9216 14522 9280
rect 14586 9216 14602 9280
rect 14666 9216 14682 9280
rect 14746 9216 14762 9280
rect 14826 9216 14834 9280
rect 14514 8192 14834 9216
rect 14514 8128 14522 8192
rect 14586 8128 14602 8192
rect 14666 8128 14682 8192
rect 14746 8128 14762 8192
rect 14826 8128 14834 8192
rect 14514 7104 14834 8128
rect 14514 7040 14522 7104
rect 14586 7040 14602 7104
rect 14666 7040 14682 7104
rect 14746 7040 14762 7104
rect 14826 7040 14834 7104
rect 14514 6016 14834 7040
rect 14514 5952 14522 6016
rect 14586 5952 14602 6016
rect 14666 5952 14682 6016
rect 14746 5952 14762 6016
rect 14826 5952 14834 6016
rect 14514 4928 14834 5952
rect 14514 4864 14522 4928
rect 14586 4864 14602 4928
rect 14666 4864 14682 4928
rect 14746 4864 14762 4928
rect 14826 4864 14834 4928
rect 14514 4742 14834 4864
rect 14514 4506 14556 4742
rect 14792 4506 14834 4742
rect 14514 3840 14834 4506
rect 14514 3776 14522 3840
rect 14586 3776 14602 3840
rect 14666 3776 14682 3840
rect 14746 3776 14762 3840
rect 14826 3776 14834 3840
rect 14514 2752 14834 3776
rect 14514 2688 14522 2752
rect 14586 2688 14602 2752
rect 14666 2688 14682 2752
rect 14746 2688 14762 2752
rect 14826 2688 14834 2752
rect 14514 2128 14834 2688
rect 15174 21792 15494 21808
rect 15174 21728 15182 21792
rect 15246 21728 15262 21792
rect 15326 21728 15342 21792
rect 15406 21728 15422 21792
rect 15486 21728 15494 21792
rect 15174 20704 15494 21728
rect 15174 20640 15182 20704
rect 15246 20640 15262 20704
rect 15326 20640 15342 20704
rect 15406 20640 15422 20704
rect 15486 20640 15494 20704
rect 15174 20090 15494 20640
rect 15174 19854 15216 20090
rect 15452 19854 15494 20090
rect 15174 19616 15494 19854
rect 15174 19552 15182 19616
rect 15246 19552 15262 19616
rect 15326 19552 15342 19616
rect 15406 19552 15422 19616
rect 15486 19552 15494 19616
rect 15174 18528 15494 19552
rect 15174 18464 15182 18528
rect 15246 18464 15262 18528
rect 15326 18464 15342 18528
rect 15406 18464 15422 18528
rect 15486 18464 15494 18528
rect 15174 17440 15494 18464
rect 15174 17376 15182 17440
rect 15246 17376 15262 17440
rect 15326 17376 15342 17440
rect 15406 17376 15422 17440
rect 15486 17376 15494 17440
rect 15174 16352 15494 17376
rect 15174 16288 15182 16352
rect 15246 16288 15262 16352
rect 15326 16288 15342 16352
rect 15406 16288 15422 16352
rect 15486 16288 15494 16352
rect 15174 15264 15494 16288
rect 15174 15200 15182 15264
rect 15246 15200 15262 15264
rect 15326 15200 15342 15264
rect 15406 15200 15422 15264
rect 15486 15200 15494 15264
rect 15174 15194 15494 15200
rect 15174 14958 15216 15194
rect 15452 14958 15494 15194
rect 15174 14176 15494 14958
rect 15174 14112 15182 14176
rect 15246 14112 15262 14176
rect 15326 14112 15342 14176
rect 15406 14112 15422 14176
rect 15486 14112 15494 14176
rect 15174 13088 15494 14112
rect 15174 13024 15182 13088
rect 15246 13024 15262 13088
rect 15326 13024 15342 13088
rect 15406 13024 15422 13088
rect 15486 13024 15494 13088
rect 15174 12000 15494 13024
rect 15174 11936 15182 12000
rect 15246 11936 15262 12000
rect 15326 11936 15342 12000
rect 15406 11936 15422 12000
rect 15486 11936 15494 12000
rect 15174 10912 15494 11936
rect 15174 10848 15182 10912
rect 15246 10848 15262 10912
rect 15326 10848 15342 10912
rect 15406 10848 15422 10912
rect 15486 10848 15494 10912
rect 15174 10298 15494 10848
rect 15174 10062 15216 10298
rect 15452 10062 15494 10298
rect 15174 9824 15494 10062
rect 15174 9760 15182 9824
rect 15246 9760 15262 9824
rect 15326 9760 15342 9824
rect 15406 9760 15422 9824
rect 15486 9760 15494 9824
rect 15174 8736 15494 9760
rect 15174 8672 15182 8736
rect 15246 8672 15262 8736
rect 15326 8672 15342 8736
rect 15406 8672 15422 8736
rect 15486 8672 15494 8736
rect 15174 7648 15494 8672
rect 15174 7584 15182 7648
rect 15246 7584 15262 7648
rect 15326 7584 15342 7648
rect 15406 7584 15422 7648
rect 15486 7584 15494 7648
rect 15174 6560 15494 7584
rect 15174 6496 15182 6560
rect 15246 6496 15262 6560
rect 15326 6496 15342 6560
rect 15406 6496 15422 6560
rect 15486 6496 15494 6560
rect 15174 5472 15494 6496
rect 15174 5408 15182 5472
rect 15246 5408 15262 5472
rect 15326 5408 15342 5472
rect 15406 5408 15422 5472
rect 15486 5408 15494 5472
rect 15174 5402 15494 5408
rect 15174 5166 15216 5402
rect 15452 5166 15494 5402
rect 15174 4384 15494 5166
rect 15174 4320 15182 4384
rect 15246 4320 15262 4384
rect 15326 4320 15342 4384
rect 15406 4320 15422 4384
rect 15486 4320 15494 4384
rect 15174 3296 15494 4320
rect 15174 3232 15182 3296
rect 15246 3232 15262 3296
rect 15326 3232 15342 3296
rect 15406 3232 15422 3296
rect 15486 3232 15494 3296
rect 15174 2208 15494 3232
rect 15174 2144 15182 2208
rect 15246 2144 15262 2208
rect 15326 2144 15342 2208
rect 15406 2144 15422 2208
rect 15486 2144 15494 2208
rect 15174 2128 15494 2144
rect 19942 21248 20262 21808
rect 19942 21184 19950 21248
rect 20014 21184 20030 21248
rect 20094 21184 20110 21248
rect 20174 21184 20190 21248
rect 20254 21184 20262 21248
rect 19942 20160 20262 21184
rect 19942 20096 19950 20160
rect 20014 20096 20030 20160
rect 20094 20096 20110 20160
rect 20174 20096 20190 20160
rect 20254 20096 20262 20160
rect 19942 19430 20262 20096
rect 19942 19194 19984 19430
rect 20220 19194 20262 19430
rect 19942 19072 20262 19194
rect 19942 19008 19950 19072
rect 20014 19008 20030 19072
rect 20094 19008 20110 19072
rect 20174 19008 20190 19072
rect 20254 19008 20262 19072
rect 19942 17984 20262 19008
rect 19942 17920 19950 17984
rect 20014 17920 20030 17984
rect 20094 17920 20110 17984
rect 20174 17920 20190 17984
rect 20254 17920 20262 17984
rect 19942 16896 20262 17920
rect 19942 16832 19950 16896
rect 20014 16832 20030 16896
rect 20094 16832 20110 16896
rect 20174 16832 20190 16896
rect 20254 16832 20262 16896
rect 19942 15808 20262 16832
rect 19942 15744 19950 15808
rect 20014 15744 20030 15808
rect 20094 15744 20110 15808
rect 20174 15744 20190 15808
rect 20254 15744 20262 15808
rect 19942 14720 20262 15744
rect 19942 14656 19950 14720
rect 20014 14656 20030 14720
rect 20094 14656 20110 14720
rect 20174 14656 20190 14720
rect 20254 14656 20262 14720
rect 19942 14534 20262 14656
rect 19942 14298 19984 14534
rect 20220 14298 20262 14534
rect 19942 13632 20262 14298
rect 19942 13568 19950 13632
rect 20014 13568 20030 13632
rect 20094 13568 20110 13632
rect 20174 13568 20190 13632
rect 20254 13568 20262 13632
rect 19942 12544 20262 13568
rect 19942 12480 19950 12544
rect 20014 12480 20030 12544
rect 20094 12480 20110 12544
rect 20174 12480 20190 12544
rect 20254 12480 20262 12544
rect 19942 11456 20262 12480
rect 19942 11392 19950 11456
rect 20014 11392 20030 11456
rect 20094 11392 20110 11456
rect 20174 11392 20190 11456
rect 20254 11392 20262 11456
rect 19942 10368 20262 11392
rect 19942 10304 19950 10368
rect 20014 10304 20030 10368
rect 20094 10304 20110 10368
rect 20174 10304 20190 10368
rect 20254 10304 20262 10368
rect 19942 9638 20262 10304
rect 19942 9402 19984 9638
rect 20220 9402 20262 9638
rect 19942 9280 20262 9402
rect 19942 9216 19950 9280
rect 20014 9216 20030 9280
rect 20094 9216 20110 9280
rect 20174 9216 20190 9280
rect 20254 9216 20262 9280
rect 19942 8192 20262 9216
rect 19942 8128 19950 8192
rect 20014 8128 20030 8192
rect 20094 8128 20110 8192
rect 20174 8128 20190 8192
rect 20254 8128 20262 8192
rect 19942 7104 20262 8128
rect 19942 7040 19950 7104
rect 20014 7040 20030 7104
rect 20094 7040 20110 7104
rect 20174 7040 20190 7104
rect 20254 7040 20262 7104
rect 19942 6016 20262 7040
rect 19942 5952 19950 6016
rect 20014 5952 20030 6016
rect 20094 5952 20110 6016
rect 20174 5952 20190 6016
rect 20254 5952 20262 6016
rect 19942 4928 20262 5952
rect 19942 4864 19950 4928
rect 20014 4864 20030 4928
rect 20094 4864 20110 4928
rect 20174 4864 20190 4928
rect 20254 4864 20262 4928
rect 19942 4742 20262 4864
rect 19942 4506 19984 4742
rect 20220 4506 20262 4742
rect 19942 3840 20262 4506
rect 19942 3776 19950 3840
rect 20014 3776 20030 3840
rect 20094 3776 20110 3840
rect 20174 3776 20190 3840
rect 20254 3776 20262 3840
rect 19942 2752 20262 3776
rect 19942 2688 19950 2752
rect 20014 2688 20030 2752
rect 20094 2688 20110 2752
rect 20174 2688 20190 2752
rect 20254 2688 20262 2752
rect 19942 2128 20262 2688
rect 20602 21792 20922 21808
rect 20602 21728 20610 21792
rect 20674 21728 20690 21792
rect 20754 21728 20770 21792
rect 20834 21728 20850 21792
rect 20914 21728 20922 21792
rect 20602 20704 20922 21728
rect 20602 20640 20610 20704
rect 20674 20640 20690 20704
rect 20754 20640 20770 20704
rect 20834 20640 20850 20704
rect 20914 20640 20922 20704
rect 20602 20090 20922 20640
rect 20602 19854 20644 20090
rect 20880 19854 20922 20090
rect 20602 19616 20922 19854
rect 20602 19552 20610 19616
rect 20674 19552 20690 19616
rect 20754 19552 20770 19616
rect 20834 19552 20850 19616
rect 20914 19552 20922 19616
rect 20602 18528 20922 19552
rect 20602 18464 20610 18528
rect 20674 18464 20690 18528
rect 20754 18464 20770 18528
rect 20834 18464 20850 18528
rect 20914 18464 20922 18528
rect 20602 17440 20922 18464
rect 20602 17376 20610 17440
rect 20674 17376 20690 17440
rect 20754 17376 20770 17440
rect 20834 17376 20850 17440
rect 20914 17376 20922 17440
rect 20602 16352 20922 17376
rect 20602 16288 20610 16352
rect 20674 16288 20690 16352
rect 20754 16288 20770 16352
rect 20834 16288 20850 16352
rect 20914 16288 20922 16352
rect 20602 15264 20922 16288
rect 20602 15200 20610 15264
rect 20674 15200 20690 15264
rect 20754 15200 20770 15264
rect 20834 15200 20850 15264
rect 20914 15200 20922 15264
rect 20602 15194 20922 15200
rect 20602 14958 20644 15194
rect 20880 14958 20922 15194
rect 20602 14176 20922 14958
rect 20602 14112 20610 14176
rect 20674 14112 20690 14176
rect 20754 14112 20770 14176
rect 20834 14112 20850 14176
rect 20914 14112 20922 14176
rect 20602 13088 20922 14112
rect 20602 13024 20610 13088
rect 20674 13024 20690 13088
rect 20754 13024 20770 13088
rect 20834 13024 20850 13088
rect 20914 13024 20922 13088
rect 20602 12000 20922 13024
rect 20602 11936 20610 12000
rect 20674 11936 20690 12000
rect 20754 11936 20770 12000
rect 20834 11936 20850 12000
rect 20914 11936 20922 12000
rect 20602 10912 20922 11936
rect 20602 10848 20610 10912
rect 20674 10848 20690 10912
rect 20754 10848 20770 10912
rect 20834 10848 20850 10912
rect 20914 10848 20922 10912
rect 20602 10298 20922 10848
rect 20602 10062 20644 10298
rect 20880 10062 20922 10298
rect 20602 9824 20922 10062
rect 20602 9760 20610 9824
rect 20674 9760 20690 9824
rect 20754 9760 20770 9824
rect 20834 9760 20850 9824
rect 20914 9760 20922 9824
rect 20602 8736 20922 9760
rect 20602 8672 20610 8736
rect 20674 8672 20690 8736
rect 20754 8672 20770 8736
rect 20834 8672 20850 8736
rect 20914 8672 20922 8736
rect 20602 7648 20922 8672
rect 20602 7584 20610 7648
rect 20674 7584 20690 7648
rect 20754 7584 20770 7648
rect 20834 7584 20850 7648
rect 20914 7584 20922 7648
rect 20602 6560 20922 7584
rect 20602 6496 20610 6560
rect 20674 6496 20690 6560
rect 20754 6496 20770 6560
rect 20834 6496 20850 6560
rect 20914 6496 20922 6560
rect 20602 5472 20922 6496
rect 20602 5408 20610 5472
rect 20674 5408 20690 5472
rect 20754 5408 20770 5472
rect 20834 5408 20850 5472
rect 20914 5408 20922 5472
rect 20602 5402 20922 5408
rect 20602 5166 20644 5402
rect 20880 5166 20922 5402
rect 20602 4384 20922 5166
rect 20602 4320 20610 4384
rect 20674 4320 20690 4384
rect 20754 4320 20770 4384
rect 20834 4320 20850 4384
rect 20914 4320 20922 4384
rect 20602 3296 20922 4320
rect 20602 3232 20610 3296
rect 20674 3232 20690 3296
rect 20754 3232 20770 3296
rect 20834 3232 20850 3296
rect 20914 3232 20922 3296
rect 20602 2208 20922 3232
rect 20602 2144 20610 2208
rect 20674 2144 20690 2208
rect 20754 2144 20770 2208
rect 20834 2144 20850 2208
rect 20914 2144 20922 2208
rect 20602 2128 20922 2144
<< via4 >>
rect 3700 19194 3936 19430
rect 3700 14298 3936 14534
rect 3700 9402 3936 9638
rect 3700 4506 3936 4742
rect 4360 19854 4596 20090
rect 4360 14958 4596 15194
rect 4360 10062 4596 10298
rect 4360 5166 4596 5402
rect 9128 19194 9364 19430
rect 9128 14298 9364 14534
rect 9128 9402 9364 9638
rect 9128 4506 9364 4742
rect 9788 19854 10024 20090
rect 9788 14958 10024 15194
rect 9788 10062 10024 10298
rect 9788 5166 10024 5402
rect 14556 19194 14792 19430
rect 14556 14298 14792 14534
rect 14556 9402 14792 9638
rect 14556 4506 14792 4742
rect 15216 19854 15452 20090
rect 15216 14958 15452 15194
rect 15216 10062 15452 10298
rect 15216 5166 15452 5402
rect 19984 19194 20220 19430
rect 19984 14298 20220 14534
rect 19984 9402 20220 9638
rect 19984 4506 20220 4742
rect 20644 19854 20880 20090
rect 20644 14958 20880 15194
rect 20644 10062 20880 10298
rect 20644 5166 20880 5402
<< metal5 >>
rect 1056 20090 22864 20132
rect 1056 19854 4360 20090
rect 4596 19854 9788 20090
rect 10024 19854 15216 20090
rect 15452 19854 20644 20090
rect 20880 19854 22864 20090
rect 1056 19812 22864 19854
rect 1056 19430 22864 19472
rect 1056 19194 3700 19430
rect 3936 19194 9128 19430
rect 9364 19194 14556 19430
rect 14792 19194 19984 19430
rect 20220 19194 22864 19430
rect 1056 19152 22864 19194
rect 1056 15194 22864 15236
rect 1056 14958 4360 15194
rect 4596 14958 9788 15194
rect 10024 14958 15216 15194
rect 15452 14958 20644 15194
rect 20880 14958 22864 15194
rect 1056 14916 22864 14958
rect 1056 14534 22864 14576
rect 1056 14298 3700 14534
rect 3936 14298 9128 14534
rect 9364 14298 14556 14534
rect 14792 14298 19984 14534
rect 20220 14298 22864 14534
rect 1056 14256 22864 14298
rect 1056 10298 22864 10340
rect 1056 10062 4360 10298
rect 4596 10062 9788 10298
rect 10024 10062 15216 10298
rect 15452 10062 20644 10298
rect 20880 10062 22864 10298
rect 1056 10020 22864 10062
rect 1056 9638 22864 9680
rect 1056 9402 3700 9638
rect 3936 9402 9128 9638
rect 9364 9402 14556 9638
rect 14792 9402 19984 9638
rect 20220 9402 22864 9638
rect 1056 9360 22864 9402
rect 1056 5402 22864 5444
rect 1056 5166 4360 5402
rect 4596 5166 9788 5402
rect 10024 5166 15216 5402
rect 15452 5166 20644 5402
rect 20880 5166 22864 5402
rect 1056 5124 22864 5166
rect 1056 4742 22864 4784
rect 1056 4506 3700 4742
rect 3936 4506 9128 4742
rect 9364 4506 14556 4742
rect 14792 4506 19984 4742
rect 20220 4506 22864 4742
rect 1056 4464 22864 4506
use sky130_fd_sc_hd__nor3b_1  _04_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 17204 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_1  _05_
timestamp 1723858470
transform 1 0 3864 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _06_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 17756 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _07_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 19228 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_1  _08_
timestamp 1723858470
transform -1 0 8556 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _09_
timestamp 1723858470
transform -1 0 4876 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _10_
timestamp 1723858470
transform 1 0 4232 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _11_
timestamp 1723858470
transform 1 0 10304 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _12_
timestamp 1723858470
transform -1 0 11040 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _13_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 17940 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _14_
timestamp 1723858470
transform -1 0 19136 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _15_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 17664 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 1932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1723858470
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1723858470
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1723858470
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1723858470
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1723858470
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_91
timestamp 1723858470
transform 1 0 9476 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_103 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 10580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 1723858470
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1723858470
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1723858470
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1723858470
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1723858470
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1723858470
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1723858470
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_169 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_177
timestamp 1723858470
transform 1 0 17388 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_189
timestamp 1723858470
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_195
timestamp 1723858470
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1723858470
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1723858470
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1723858470
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_225
timestamp 1723858470
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1723858470
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1723858470
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1723858470
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1723858470
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1723858470
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1723858470
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1723858470
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1723858470
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1723858470
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1723858470
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1723858470
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1723858470
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1723858470
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1723858470
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1723858470
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1723858470
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1723858470
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1723858470
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1723858470
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1723858470
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1723858470
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1723858470
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1723858470
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_225
timestamp 1723858470
transform 1 0 21804 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1723858470
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1723858470
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1723858470
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1723858470
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1723858470
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1723858470
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1723858470
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1723858470
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1723858470
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1723858470
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1723858470
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1723858470
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1723858470
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1723858470
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1723858470
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1723858470
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1723858470
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1723858470
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1723858470
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1723858470
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1723858470
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1723858470
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1723858470
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1723858470
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1723858470
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1723858470
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1723858470
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1723858470
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1723858470
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1723858470
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1723858470
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_69
timestamp 1723858470
transform 1 0 7452 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1723858470
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1723858470
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1723858470
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1723858470
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1723858470
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1723858470
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1723858470
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1723858470
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1723858470
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1723858470
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1723858470
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1723858470
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1723858470
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1723858470
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1723858470
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1723858470
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_225
timestamp 1723858470
transform 1 0 21804 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1723858470
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1723858470
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1723858470
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1723858470
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1723858470
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1723858470
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1723858470
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1723858470
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1723858470
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1723858470
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1723858470
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1723858470
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1723858470
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1723858470
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1723858470
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1723858470
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1723858470
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1723858470
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1723858470
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1723858470
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1723858470
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1723858470
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1723858470
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1723858470
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1723858470
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1723858470
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1723858470
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1723858470
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1723858470
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1723858470
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1723858470
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1723858470
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1723858470
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1723858470
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1723858470
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1723858470
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1723858470
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1723858470
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1723858470
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1723858470
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1723858470
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1723858470
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_175
timestamp 1723858470
transform 1 0 17204 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_187
timestamp 1723858470
transform 1 0 18308 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_199
timestamp 1723858470
transform 1 0 19412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_211
timestamp 1723858470
transform 1 0 20516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1723858470
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_225
timestamp 1723858470
transform 1 0 21804 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1723858470
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1723858470
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1723858470
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1723858470
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1723858470
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1723858470
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1723858470
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1723858470
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1723858470
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1723858470
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1723858470
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1723858470
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1723858470
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1723858470
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1723858470
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1723858470
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1723858470
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1723858470
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1723858470
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1723858470
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1723858470
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1723858470
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1723858470
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1723858470
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1723858470
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1723858470
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1723858470
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1723858470
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1723858470
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1723858470
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1723858470
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1723858470
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1723858470
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1723858470
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1723858470
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1723858470
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1723858470
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1723858470
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1723858470
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1723858470
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1723858470
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1723858470
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1723858470
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1723858470
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1723858470
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1723858470
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1723858470
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1723858470
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_225
timestamp 1723858470
transform 1 0 21804 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1723858470
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1723858470
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1723858470
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1723858470
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1723858470
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1723858470
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1723858470
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1723858470
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1723858470
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1723858470
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1723858470
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1723858470
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1723858470
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1723858470
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1723858470
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1723858470
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1723858470
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1723858470
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1723858470
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1723858470
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1723858470
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1723858470
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1723858470
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1723858470
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1723858470
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1723858470
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1723858470
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1723858470
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1723858470
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1723858470
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1723858470
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1723858470
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1723858470
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1723858470
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1723858470
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1723858470
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1723858470
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1723858470
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1723858470
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1723858470
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1723858470
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1723858470
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1723858470
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1723858470
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1723858470
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1723858470
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1723858470
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1723858470
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_225
timestamp 1723858470
transform 1 0 21804 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1723858470
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1723858470
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1723858470
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1723858470
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1723858470
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1723858470
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1723858470
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1723858470
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1723858470
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1723858470
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1723858470
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1723858470
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1723858470
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1723858470
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1723858470
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1723858470
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1723858470
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1723858470
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1723858470
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1723858470
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1723858470
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1723858470
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1723858470
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1723858470
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1723858470
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1723858470
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1723858470
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1723858470
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1723858470
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1723858470
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1723858470
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1723858470
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1723858470
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1723858470
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1723858470
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1723858470
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1723858470
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1723858470
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1723858470
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1723858470
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1723858470
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1723858470
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1723858470
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1723858470
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1723858470
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1723858470
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1723858470
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1723858470
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_225
timestamp 1723858470
transform 1 0 21804 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_9
timestamp 1723858470
transform 1 0 1932 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_21
timestamp 1723858470
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1723858470
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_29
timestamp 1723858470
transform 1 0 3772 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_36
timestamp 1723858470
transform 1 0 4416 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_48
timestamp 1723858470
transform 1 0 5520 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_60
timestamp 1723858470
transform 1 0 6624 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_72
timestamp 1723858470
transform 1 0 7728 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1723858470
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1723858470
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1723858470
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1723858470
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1723858470
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1723858470
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1723858470
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1723858470
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1723858470
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1723858470
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1723858470
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1723858470
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1723858470
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 1723858470
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 1723858470
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1723858470
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1723858470
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1723858470
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1723858470
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1723858470
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1723858470
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1723858470
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1723858470
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1723858470
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1723858470
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1723858470
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1723858470
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1723858470
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1723858470
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 1723858470
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_149
timestamp 1723858470
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_161
timestamp 1723858470
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1723858470
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1723858470
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_181
timestamp 1723858470
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_193
timestamp 1723858470
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_205
timestamp 1723858470
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_217
timestamp 1723858470
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1723858470
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_225
timestamp 1723858470
transform 1 0 21804 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1723858470
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1723858470
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1723858470
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1723858470
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1723858470
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1723858470
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1723858470
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1723858470
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1723858470
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1723858470
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1723858470
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1723858470
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1723858470
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1723858470
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1723858470
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1723858470
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 1723858470
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 1723858470
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_177
timestamp 1723858470
transform 1 0 17388 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_188
timestamp 1723858470
transform 1 0 18400 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 1723858470
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_209
timestamp 1723858470
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_221
timestamp 1723858470
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1723858470
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1723858470
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1723858470
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1723858470
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1723858470
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1723858470
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1723858470
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1723858470
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1723858470
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 1723858470
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1723858470
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1723858470
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1723858470
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1723858470
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 1723858470
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 1723858470
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_161
timestamp 1723858470
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1723858470
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 1723858470
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_181
timestamp 1723858470
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_196
timestamp 1723858470
transform 1 0 19136 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_208
timestamp 1723858470
transform 1 0 20240 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_220
timestamp 1723858470
transform 1 0 21344 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_225
timestamp 1723858470
transform 1 0 21804 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1723858470
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1723858470
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1723858470
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1723858470
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1723858470
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1723858470
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1723858470
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1723858470
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1723858470
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1723858470
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1723858470
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 1723858470
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 1723858470
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 1723858470
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1723858470
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 1723858470
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_153
timestamp 1723858470
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_165
timestamp 1723858470
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_177
timestamp 1723858470
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_189
timestamp 1723858470
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1723858470
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_197
timestamp 1723858470
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_209
timestamp 1723858470
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_221
timestamp 1723858470
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1723858470
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1723858470
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1723858470
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1723858470
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1723858470
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1723858470
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1723858470
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1723858470
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1723858470
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1723858470
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 1723858470
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1723858470
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1723858470
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 1723858470
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_137
timestamp 1723858470
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_149
timestamp 1723858470
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_161
timestamp 1723858470
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1723858470
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1723858470
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_181
timestamp 1723858470
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_193
timestamp 1723858470
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_205
timestamp 1723858470
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_217
timestamp 1723858470
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 1723858470
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_225
timestamp 1723858470
transform 1 0 21804 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1723858470
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1723858470
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1723858470
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1723858470
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1723858470
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1723858470
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1723858470
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 1723858470
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1723858470
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1723858470
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1723858470
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 1723858470
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_121
timestamp 1723858470
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 1723858470
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1723858470
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1723858470
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_153
timestamp 1723858470
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_165
timestamp 1723858470
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_177
timestamp 1723858470
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_189
timestamp 1723858470
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 1723858470
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_197
timestamp 1723858470
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_209
timestamp 1723858470
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_221
timestamp 1723858470
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1723858470
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1723858470
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1723858470
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1723858470
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1723858470
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1723858470
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1723858470
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1723858470
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 1723858470
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 1723858470
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 1723858470
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1723858470
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 1723858470
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 1723858470
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_137
timestamp 1723858470
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_149
timestamp 1723858470
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_161
timestamp 1723858470
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1723858470
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 1723858470
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_181
timestamp 1723858470
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_193
timestamp 1723858470
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_205
timestamp 1723858470
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_217
timestamp 1723858470
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 1723858470
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_225
timestamp 1723858470
transform 1 0 21804 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1723858470
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1723858470
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1723858470
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1723858470
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1723858470
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1723858470
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1723858470
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1723858470
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1723858470
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1723858470
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 1723858470
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_109
timestamp 1723858470
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_121
timestamp 1723858470
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_133
timestamp 1723858470
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1723858470
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1723858470
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_153
timestamp 1723858470
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_165
timestamp 1723858470
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_177
timestamp 1723858470
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_189
timestamp 1723858470
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1723858470
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_197
timestamp 1723858470
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_209
timestamp 1723858470
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_221
timestamp 1723858470
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1723858470
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1723858470
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1723858470
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1723858470
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1723858470
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1723858470
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1723858470
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1723858470
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 1723858470
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 1723858470
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 1723858470
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1723858470
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1723858470
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 1723858470
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_137
timestamp 1723858470
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_149
timestamp 1723858470
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_161
timestamp 1723858470
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1723858470
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1723858470
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_181
timestamp 1723858470
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_193
timestamp 1723858470
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_205
timestamp 1723858470
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_217
timestamp 1723858470
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1723858470
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_225
timestamp 1723858470
transform 1 0 21804 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1723858470
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1723858470
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1723858470
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1723858470
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1723858470
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1723858470
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 1723858470
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 1723858470
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1723858470
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1723858470
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 1723858470
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_109
timestamp 1723858470
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_121
timestamp 1723858470
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_133
timestamp 1723858470
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1723858470
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1723858470
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_153
timestamp 1723858470
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_165
timestamp 1723858470
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_177
timestamp 1723858470
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_189
timestamp 1723858470
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1723858470
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_197
timestamp 1723858470
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_209
timestamp 1723858470
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_221
timestamp 1723858470
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1723858470
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1723858470
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1723858470
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1723858470
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1723858470
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1723858470
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1723858470
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1723858470
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 1723858470
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 1723858470
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 1723858470
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1723858470
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1723858470
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 1723858470
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_137
timestamp 1723858470
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_149
timestamp 1723858470
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 1723858470
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1723858470
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 1723858470
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_181
timestamp 1723858470
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_193
timestamp 1723858470
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_205
timestamp 1723858470
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_217
timestamp 1723858470
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1723858470
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_225
timestamp 1723858470
transform 1 0 21804 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1723858470
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1723858470
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1723858470
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1723858470
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1723858470
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 1723858470
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 1723858470
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 1723858470
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1723858470
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1723858470
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 1723858470
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_109
timestamp 1723858470
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_121
timestamp 1723858470
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 1723858470
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1723858470
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 1723858470
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_153
timestamp 1723858470
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_165
timestamp 1723858470
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_177
timestamp 1723858470
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_189
timestamp 1723858470
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 1723858470
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 1723858470
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_209
timestamp 1723858470
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_221
timestamp 1723858470
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1723858470
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1723858470
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1723858470
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1723858470
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1723858470
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1723858470
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1723858470
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1723858470
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1723858470
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 1723858470
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 1723858470
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1723858470
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1723858470
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 1723858470
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_137
timestamp 1723858470
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 1723858470
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 1723858470
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1723858470
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1723858470
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp 1723858470
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_193
timestamp 1723858470
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_205
timestamp 1723858470
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_217
timestamp 1723858470
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1723858470
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_225
timestamp 1723858470
transform 1 0 21804 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1723858470
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1723858470
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1723858470
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1723858470
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1723858470
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1723858470
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1723858470
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 1723858470
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1723858470
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1723858470
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 1723858470
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 1723858470
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 1723858470
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 1723858470
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1723858470
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1723858470
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 1723858470
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 1723858470
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_177
timestamp 1723858470
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_189
timestamp 1723858470
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 1723858470
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 1723858470
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_209
timestamp 1723858470
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_221
timestamp 1723858470
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1723858470
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1723858470
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 1723858470
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 1723858470
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 1723858470
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1723858470
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1723858470
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1723858470
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_81
timestamp 1723858470
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_93
timestamp 1723858470
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_105
timestamp 1723858470
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1723858470
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 1723858470
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 1723858470
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_137
timestamp 1723858470
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_149
timestamp 1723858470
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_161
timestamp 1723858470
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1723858470
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1723858470
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_181
timestamp 1723858470
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_193
timestamp 1723858470
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_205
timestamp 1723858470
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_217
timestamp 1723858470
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1723858470
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_225
timestamp 1723858470
transform 1 0 21804 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1723858470
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1723858470
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1723858470
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1723858470
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1723858470
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 1723858470
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 1723858470
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 1723858470
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1723858470
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1723858470
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 1723858470
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_109
timestamp 1723858470
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_121
timestamp 1723858470
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_133
timestamp 1723858470
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1723858470
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 1723858470
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_153
timestamp 1723858470
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_165
timestamp 1723858470
transform 1 0 16284 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_173
timestamp 1723858470
transform 1 0 17020 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_180
timestamp 1723858470
transform 1 0 17664 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_188
timestamp 1723858470
transform 1 0 18400 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 1723858470
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_209
timestamp 1723858470
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_221
timestamp 1723858470
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_9
timestamp 1723858470
transform 1 0 1932 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_21
timestamp 1723858470
transform 1 0 3036 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_33
timestamp 1723858470
transform 1 0 4140 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_41
timestamp 1723858470
transform 1 0 4876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_53
timestamp 1723858470
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1723858470
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 1723858470
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_81
timestamp 1723858470
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_93
timestamp 1723858470
transform 1 0 9660 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_99
timestamp 1723858470
transform 1 0 10212 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_107
timestamp 1723858470
transform 1 0 10948 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1723858470
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1723858470
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 1723858470
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_137
timestamp 1723858470
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_149
timestamp 1723858470
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_161
timestamp 1723858470
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1723858470
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1723858470
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_181
timestamp 1723858470
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_193
timestamp 1723858470
transform 1 0 18860 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_197
timestamp 1723858470
transform 1 0 19228 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_209
timestamp 1723858470
transform 1 0 20332 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_221
timestamp 1723858470
transform 1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_225
timestamp 1723858470
transform 1 0 21804 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1723858470
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1723858470
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1723858470
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_29
timestamp 1723858470
transform 1 0 3772 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_33
timestamp 1723858470
transform 1 0 4140 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_37
timestamp 1723858470
transform 1 0 4508 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_49
timestamp 1723858470
transform 1 0 5612 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_61
timestamp 1723858470
transform 1 0 6716 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_73
timestamp 1723858470
transform 1 0 7820 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_81
timestamp 1723858470
transform 1 0 8556 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1723858470
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_97
timestamp 1723858470
transform 1 0 10028 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_108
timestamp 1723858470
transform 1 0 11040 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_120
timestamp 1723858470
transform 1 0 12144 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_132
timestamp 1723858470
transform 1 0 13248 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1723858470
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 1723858470
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_165
timestamp 1723858470
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_177
timestamp 1723858470
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_189
timestamp 1723858470
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 1723858470
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_197
timestamp 1723858470
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_209
timestamp 1723858470
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_221
timestamp 1723858470
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1723858470
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1723858470
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 1723858470
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 1723858470
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 1723858470
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1723858470
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1723858470
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 1723858470
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 1723858470
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_93
timestamp 1723858470
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_105
timestamp 1723858470
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1723858470
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 1723858470
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_125
timestamp 1723858470
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_137
timestamp 1723858470
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_149
timestamp 1723858470
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_161
timestamp 1723858470
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1723858470
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1723858470
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_181
timestamp 1723858470
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_193
timestamp 1723858470
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_205
timestamp 1723858470
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_217
timestamp 1723858470
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 1723858470
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_225
timestamp 1723858470
transform 1 0 21804 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1723858470
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1723858470
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1723858470
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1723858470
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1723858470
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 1723858470
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_65
timestamp 1723858470
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 1723858470
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1723858470
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1723858470
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_97
timestamp 1723858470
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_109
timestamp 1723858470
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_121
timestamp 1723858470
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_133
timestamp 1723858470
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1723858470
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 1723858470
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_153
timestamp 1723858470
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_165
timestamp 1723858470
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_177
timestamp 1723858470
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_189
timestamp 1723858470
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1723858470
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 1723858470
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_209
timestamp 1723858470
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_221
timestamp 1723858470
transform 1 0 21436 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1723858470
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1723858470
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 1723858470
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_39
timestamp 1723858470
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 1723858470
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1723858470
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1723858470
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1723858470
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_81
timestamp 1723858470
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_93
timestamp 1723858470
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_105
timestamp 1723858470
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1723858470
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 1723858470
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_125
timestamp 1723858470
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_137
timestamp 1723858470
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_149
timestamp 1723858470
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_161
timestamp 1723858470
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 1723858470
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 1723858470
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_181
timestamp 1723858470
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_193
timestamp 1723858470
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_205
timestamp 1723858470
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_217
timestamp 1723858470
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_223
timestamp 1723858470
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_225
timestamp 1723858470
transform 1 0 21804 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1723858470
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 1723858470
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1723858470
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 1723858470
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_41
timestamp 1723858470
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_53
timestamp 1723858470
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_65
timestamp 1723858470
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_77
timestamp 1723858470
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 1723858470
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_85
timestamp 1723858470
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_97
timestamp 1723858470
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_109
timestamp 1723858470
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_121
timestamp 1723858470
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_133
timestamp 1723858470
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 1723858470
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_141
timestamp 1723858470
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_153
timestamp 1723858470
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_165
timestamp 1723858470
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_177
timestamp 1723858470
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_189
timestamp 1723858470
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_195
timestamp 1723858470
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_197
timestamp 1723858470
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_209
timestamp 1723858470
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_221
timestamp 1723858470
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1723858470
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_21
timestamp 1723858470
transform 1 0 3036 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_27
timestamp 1723858470
transform 1 0 3588 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_29
timestamp 1723858470
transform 1 0 3772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_41
timestamp 1723858470
transform 1 0 4876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_53
timestamp 1723858470
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 1723858470
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_69
timestamp 1723858470
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_81
timestamp 1723858470
transform 1 0 8556 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_85
timestamp 1723858470
transform 1 0 8924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_97
timestamp 1723858470
transform 1 0 10028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_109
timestamp 1723858470
transform 1 0 11132 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_119
timestamp 1723858470
transform 1 0 12052 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_131
timestamp 1723858470
transform 1 0 13156 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_139
timestamp 1723858470
transform 1 0 13892 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_141
timestamp 1723858470
transform 1 0 14076 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_153
timestamp 1723858470
transform 1 0 15180 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_165
timestamp 1723858470
transform 1 0 16284 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 1723858470
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_181
timestamp 1723858470
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_193
timestamp 1723858470
transform 1 0 18860 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_197
timestamp 1723858470
transform 1 0 19228 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_205
timestamp 1723858470
transform 1 0 19964 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_210
timestamp 1723858470
transform 1 0 20424 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_222
timestamp 1723858470
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_225
timestamp 1723858470
transform 1 0 21804 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 1380 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input2
timestamp 1723858470
transform -1 0 22540 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input3
timestamp 1723858470
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 20056 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output5
timestamp 1723858470
transform 1 0 16836 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output6
timestamp 1723858470
transform -1 0 1932 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1723858470
transform 1 0 22172 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output8
timestamp 1723858470
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output9
timestamp 1723858470
transform -1 0 3036 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output10
timestamp 1723858470
transform 1 0 11500 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1723858470
transform 1 0 22172 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1723858470
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1723858470
transform -1 0 22816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1723858470
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1723858470
transform -1 0 22816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1723858470
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1723858470
transform -1 0 22816 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1723858470
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1723858470
transform -1 0 22816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1723858470
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1723858470
transform -1 0 22816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1723858470
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1723858470
transform -1 0 22816 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1723858470
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1723858470
transform -1 0 22816 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1723858470
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1723858470
transform -1 0 22816 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1723858470
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1723858470
transform -1 0 22816 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1723858470
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1723858470
transform -1 0 22816 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1723858470
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1723858470
transform -1 0 22816 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1723858470
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1723858470
transform -1 0 22816 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1723858470
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1723858470
transform -1 0 22816 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1723858470
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1723858470
transform -1 0 22816 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1723858470
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1723858470
transform -1 0 22816 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1723858470
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1723858470
transform -1 0 22816 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1723858470
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1723858470
transform -1 0 22816 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1723858470
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1723858470
transform -1 0 22816 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1723858470
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1723858470
transform -1 0 22816 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1723858470
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1723858470
transform -1 0 22816 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1723858470
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1723858470
transform -1 0 22816 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1723858470
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1723858470
transform -1 0 22816 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1723858470
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1723858470
transform -1 0 22816 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1723858470
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1723858470
transform -1 0 22816 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1723858470
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1723858470
transform -1 0 22816 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1723858470
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1723858470
transform -1 0 22816 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1723858470
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1723858470
transform -1 0 22816 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1723858470
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1723858470
transform -1 0 22816 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1723858470
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1723858470
transform -1 0 22816 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1723858470
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1723858470
transform -1 0 22816 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1723858470
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1723858470
transform -1 0 22816 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1723858470
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1723858470
transform -1 0 22816 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1723858470
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1723858470
transform -1 0 22816 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1723858470
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1723858470
transform -1 0 22816 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1723858470
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1723858470
transform -1 0 22816 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1723858470
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1723858470
transform -1 0 22816 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1723858470
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1723858470
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1723858470
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1723858470
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1723858470
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1723858470
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1723858470
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1723858470
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1723858470
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1723858470
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1723858470
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1723858470
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1723858470
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1723858470
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1723858470
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1723858470
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1723858470
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1723858470
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1723858470
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1723858470
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1723858470
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1723858470
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1723858470
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1723858470
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1723858470
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1723858470
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1723858470
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1723858470
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1723858470
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1723858470
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1723858470
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1723858470
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1723858470
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1723858470
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1723858470
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1723858470
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1723858470
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1723858470
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1723858470
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1723858470
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1723858470
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1723858470
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1723858470
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1723858470
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1723858470
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1723858470
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1723858470
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1723858470
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1723858470
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1723858470
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1723858470
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1723858470
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1723858470
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1723858470
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1723858470
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1723858470
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1723858470
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1723858470
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1723858470
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1723858470
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1723858470
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1723858470
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1723858470
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1723858470
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1723858470
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1723858470
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1723858470
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1723858470
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1723858470
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1723858470
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1723858470
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1723858470
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1723858470
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1723858470
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1723858470
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1723858470
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1723858470
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1723858470
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1723858470
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1723858470
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1723858470
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1723858470
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1723858470
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1723858470
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1723858470
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1723858470
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1723858470
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1723858470
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1723858470
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1723858470
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1723858470
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1723858470
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1723858470
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1723858470
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1723858470
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1723858470
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1723858470
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1723858470
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1723858470
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1723858470
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1723858470
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1723858470
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1723858470
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1723858470
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1723858470
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1723858470
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1723858470
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1723858470
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1723858470
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1723858470
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1723858470
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1723858470
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1723858470
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1723858470
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1723858470
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1723858470
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1723858470
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1723858470
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1723858470
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1723858470
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1723858470
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1723858470
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1723858470
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1723858470
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1723858470
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1723858470
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1723858470
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1723858470
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1723858470
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1723858470
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1723858470
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1723858470
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1723858470
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1723858470
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1723858470
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1723858470
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1723858470
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1723858470
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1723858470
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1723858470
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1723858470
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1723858470
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1723858470
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1723858470
transform 1 0 3680 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1723858470
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1723858470
transform 1 0 8832 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1723858470
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1723858470
transform 1 0 13984 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1723858470
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1723858470
transform 1 0 19136 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1723858470
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
<< labels >>
flabel metal4 s 4318 2128 4638 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 9746 2128 10066 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 15174 2128 15494 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 20602 2128 20922 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 5124 22864 5444 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 10020 22864 10340 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 14916 22864 15236 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 19812 22864 20132 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 3658 2128 3978 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 9086 2128 9406 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 14514 2128 14834 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 19942 2128 20262 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 4464 22864 4784 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 9360 22864 9680 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 14256 22864 14576 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 19152 22864 19472 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 in[0]
port 2 nsew signal input
flabel metal3 s 23200 1368 24000 1488 0 FreeSans 480 0 0 0 in[1]
port 3 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 in[2]
port 4 nsew signal input
flabel metal2 s 19982 23200 20038 24000 0 FreeSans 224 90 0 0 out[0]
port 5 nsew signal tristate
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 out[1]
port 6 nsew signal tristate
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 out[2]
port 7 nsew signal tristate
flabel metal3 s 23200 19728 24000 19848 0 FreeSans 480 0 0 0 out[3]
port 8 nsew signal tristate
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 out[4]
port 9 nsew signal tristate
flabel metal2 s 2594 23200 2650 24000 0 FreeSans 224 90 0 0 out[5]
port 10 nsew signal tristate
flabel metal2 s 10966 23200 11022 24000 0 FreeSans 224 90 0 0 out[6]
port 11 nsew signal tristate
flabel metal3 s 23200 10208 24000 10328 0 FreeSans 480 0 0 0 out[7]
port 12 nsew signal tristate
rlabel metal1 11960 21760 11960 21760 0 VGND
rlabel metal1 11960 21216 11960 21216 0 VPWR
rlabel metal1 18676 17850 18676 17850 0 _00_
rlabel metal2 4278 18564 4278 18564 0 _01_
rlabel metal1 10856 18394 10856 18394 0 _02_
rlabel metal1 18630 10234 18630 10234 0 _03_
rlabel metal3 751 17748 751 17748 0 in[0]
rlabel metal1 22632 2346 22632 2346 0 in[1]
rlabel metal2 46 1554 46 1554 0 in[2]
rlabel metal1 17526 5270 17526 5270 0 net1
rlabel metal2 10994 20230 10994 20230 0 net10
rlabel metal1 20654 10642 20654 10642 0 net11
rlabel metal2 22126 3366 22126 3366 0 net2
rlabel metal1 3266 2618 3266 2618 0 net3
rlabel metal1 17848 17850 17848 17850 0 net4
rlabel metal1 17066 2414 17066 2414 0 net5
rlabel metal1 2852 8874 2852 8874 0 net6
rlabel metal1 20700 18394 20700 18394 0 net7
rlabel metal1 8786 2414 8786 2414 0 net8
rlabel metal2 4278 20230 4278 20230 0 net9
rlabel metal2 20286 22491 20286 22491 0 out[0]
rlabel metal2 16790 1520 16790 1520 0 out[1]
rlabel metal3 820 8908 820 8908 0 out[2]
rlabel metal1 22632 20026 22632 20026 0 out[3]
rlabel metal2 8418 1520 8418 1520 0 out[4]
rlabel metal2 2622 22484 2622 22484 0 out[5]
rlabel metal2 10994 22695 10994 22695 0 out[6]
rlabel metal2 22402 10353 22402 10353 0 out[7]
<< properties >>
string FIXED_BBOX 0 0 24000 24000
<< end >>
