magic
tech sky130A
magscale 1 2
timestamp 1755279893
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 14 2128 38994 37584
<< metal2 >>
rect 3882 39200 3938 40000
rect 18050 39200 18106 40000
rect 32218 39200 32274 40000
rect 18 0 74 800
rect 14186 0 14242 800
rect 28354 0 28410 800
<< obsm2 >>
rect 20 39144 3826 39200
rect 3994 39144 17994 39200
rect 18162 39144 32162 39200
rect 32330 39144 38990 39200
rect 20 856 38990 39144
rect 130 800 14130 856
rect 14298 800 28298 856
rect 28466 800 38990 856
<< metal3 >>
rect 39200 32648 40000 32768
rect 0 29248 800 29368
rect 39200 17688 40000 17808
rect 0 14288 800 14408
rect 39200 2728 40000 2848
<< obsm3 >>
rect 800 32848 39200 37569
rect 800 32568 39120 32848
rect 800 29448 39200 32568
rect 880 29168 39200 29448
rect 800 17888 39200 29168
rect 800 17608 39120 17888
rect 800 14488 39200 17608
rect 880 14208 39200 14488
rect 800 2928 39200 14208
rect 800 2648 39120 2928
rect 800 2143 39200 2648
<< metal4 >>
rect 4208 2128 4528 37584
rect 4868 2128 5188 37584
rect 34928 2128 35248 37584
rect 35588 2128 35908 37584
<< metal5 >>
rect 1056 36642 38872 36962
rect 1056 35982 38872 36302
rect 1056 6006 38872 6326
rect 1056 5346 38872 5666
<< labels >>
rlabel metal4 s 4868 2128 5188 37584 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 35588 2128 35908 37584 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 6006 38872 6326 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 36642 38872 36962 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 37584 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 5346 38872 5666 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 35982 38872 36302 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 29248 800 29368 6 in[0]
port 3 nsew signal input
rlabel metal3 s 39200 2728 40000 2848 6 in[1]
port 4 nsew signal input
rlabel metal2 s 18 0 74 800 6 in[2]
port 5 nsew signal input
rlabel metal2 s 32218 39200 32274 40000 6 out[0]
port 6 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 out[1]
port 7 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 out[2]
port 8 nsew signal output
rlabel metal3 s 39200 32648 40000 32768 6 out[3]
port 9 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 out[4]
port 10 nsew signal output
rlabel metal2 s 3882 39200 3938 40000 6 out[5]
port 11 nsew signal output
rlabel metal2 s 18050 39200 18106 40000 6 out[6]
port 12 nsew signal output
rlabel metal3 s 39200 17688 40000 17808 6 out[7]
port 13 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 516306
string GDS_FILE /openlane/designs/decoder3to8/runs/run1//results/signoff/decoder3to8.magic.gds
string GDS_START 65868
<< end >>

