magic
tech sky130A
magscale 1 2
timestamp 1755207336
<< obsli1 >>
rect 1104 2159 22816 21777
<< obsm1 >>
rect 14 2128 22894 21808
<< metal2 >>
rect 2594 23200 2650 24000
rect 10966 23200 11022 24000
rect 19982 23200 20038 24000
rect 18 0 74 800
rect 8390 0 8446 800
rect 16762 0 16818 800
<< obsm2 >>
rect 20 23144 2538 23338
rect 2706 23144 10910 23338
rect 11078 23144 19926 23338
rect 20094 23144 22890 23338
rect 20 856 22890 23144
rect 130 800 8334 856
rect 8502 800 16706 856
rect 16874 800 22890 856
<< metal3 >>
rect 23200 19728 24000 19848
rect 0 17688 800 17808
rect 23200 10208 24000 10328
rect 0 8848 800 8968
rect 23200 1368 24000 1488
<< obsm3 >>
rect 798 19928 23200 21793
rect 798 19648 23120 19928
rect 798 17888 23200 19648
rect 880 17608 23200 17888
rect 798 10408 23200 17608
rect 798 10128 23120 10408
rect 798 9048 23200 10128
rect 880 8768 23200 9048
rect 798 1568 23200 8768
rect 798 1395 23120 1568
<< metal4 >>
rect 3658 2128 3978 21808
rect 4318 2128 4638 21808
rect 9086 2128 9406 21808
rect 9746 2128 10066 21808
rect 14514 2128 14834 21808
rect 15174 2128 15494 21808
rect 19942 2128 20262 21808
rect 20602 2128 20922 21808
<< metal5 >>
rect 1056 19812 22864 20132
rect 1056 19152 22864 19472
rect 1056 14916 22864 15236
rect 1056 14256 22864 14576
rect 1056 10020 22864 10340
rect 1056 9360 22864 9680
rect 1056 5124 22864 5444
rect 1056 4464 22864 4784
<< labels >>
rlabel metal4 s 4318 2128 4638 21808 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 9746 2128 10066 21808 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 15174 2128 15494 21808 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 20602 2128 20922 21808 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 5124 22864 5444 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 10020 22864 10340 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 14916 22864 15236 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 19812 22864 20132 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 3658 2128 3978 21808 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 9086 2128 9406 21808 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 14514 2128 14834 21808 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 19942 2128 20262 21808 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 4464 22864 4784 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 9360 22864 9680 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 14256 22864 14576 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 19152 22864 19472 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 17688 800 17808 6 in[0]
port 3 nsew signal input
rlabel metal3 s 23200 1368 24000 1488 6 in[1]
port 4 nsew signal input
rlabel metal2 s 18 0 74 800 6 in[2]
port 5 nsew signal input
rlabel metal2 s 19982 23200 20038 24000 6 out[0]
port 6 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 out[1]
port 7 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 out[2]
port 8 nsew signal output
rlabel metal3 s 23200 19728 24000 19848 6 out[3]
port 9 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 out[4]
port 10 nsew signal output
rlabel metal2 s 2594 23200 2650 24000 6 out[5]
port 11 nsew signal output
rlabel metal2 s 10966 23200 11022 24000 6 out[6]
port 12 nsew signal output
rlabel metal3 s 23200 10208 24000 10328 6 out[7]
port 13 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 24000 24000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 334758
string GDS_FILE /openlane/designs/decoder3to8/runs/RUN_2025.08.14_21.34.53/results/signoff/decoder3to8.magic.gds
string GDS_START 56504
<< end >>

